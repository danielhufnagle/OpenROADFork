module gcd (clk,
    req_rdy,
    req_val,
    reset,
    resp_rdy,
    resp_val,
    req_msg,
    resp_msg,
    VSS,
    VDD);
 input clk;
 output req_rdy;
 input req_val;
 input reset;
 input resp_rdy;
 output resp_val;
 input [31:0] req_msg;
 output [15:0] resp_msg;
 inout VSS;
 inout VDD;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire \ctrl.state.out[1] ;
 wire \ctrl.state.out[2] ;
 wire \dpath.a_lt_b$in0[0] ;
 wire \dpath.a_lt_b$in0[10] ;
 wire \dpath.a_lt_b$in0[11] ;
 wire \dpath.a_lt_b$in0[12] ;
 wire \dpath.a_lt_b$in0[13] ;
 wire \dpath.a_lt_b$in0[14] ;
 wire \dpath.a_lt_b$in0[15] ;
 wire \dpath.a_lt_b$in0[1] ;
 wire \dpath.a_lt_b$in0[2] ;
 wire \dpath.a_lt_b$in0[3] ;
 wire \dpath.a_lt_b$in0[4] ;
 wire \dpath.a_lt_b$in0[5] ;
 wire \dpath.a_lt_b$in0[6] ;
 wire \dpath.a_lt_b$in0[7] ;
 wire \dpath.a_lt_b$in0[8] ;
 wire \dpath.a_lt_b$in0[9] ;
 wire \dpath.a_lt_b$in1[0] ;
 wire \dpath.a_lt_b$in1[10] ;
 wire \dpath.a_lt_b$in1[11] ;
 wire \dpath.a_lt_b$in1[12] ;
 wire \dpath.a_lt_b$in1[13] ;
 wire \dpath.a_lt_b$in1[14] ;
 wire \dpath.a_lt_b$in1[15] ;
 wire \dpath.a_lt_b$in1[1] ;
 wire \dpath.a_lt_b$in1[2] ;
 wire \dpath.a_lt_b$in1[3] ;
 wire \dpath.a_lt_b$in1[4] ;
 wire \dpath.a_lt_b$in1[5] ;
 wire \dpath.a_lt_b$in1[6] ;
 wire \dpath.a_lt_b$in1[7] ;
 wire \dpath.a_lt_b$in1[8] ;
 wire \dpath.a_lt_b$in1[9] ;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 INV_X4 _345_ (.A(\dpath.a_lt_b$in1[1] ),
    .ZN(_036_));
 BUF_X4 _346_ (.A(\dpath.a_lt_b$in0[1] ),
    .Z(_037_));
 NAND2_X1 _347_ (.A1(_036_),
    .A2(_037_),
    .ZN(_038_));
 INV_X2 _348_ (.A(\dpath.a_lt_b$in1[0] ),
    .ZN(_039_));
 NOR2_X2 _349_ (.A1(_039_),
    .A2(\dpath.a_lt_b$in0[0] ),
    .ZN(_040_));
 NOR2_X2 _350_ (.A1(_036_),
    .A2(_037_),
    .ZN(_041_));
 OAI21_X4 _351_ (.A(_038_),
    .B1(_040_),
    .B2(_041_),
    .ZN(_042_));
 INV_X2 _352_ (.A(\dpath.a_lt_b$in1[3] ),
    .ZN(_043_));
 NAND2_X2 _353_ (.A1(_043_),
    .A2(\dpath.a_lt_b$in0[3] ),
    .ZN(_044_));
 INV_X2 _354_ (.A(\dpath.a_lt_b$in0[3] ),
    .ZN(_045_));
 NAND2_X2 _355_ (.A1(_045_),
    .A2(\dpath.a_lt_b$in1[3] ),
    .ZN(_046_));
 NAND2_X4 _356_ (.A1(_046_),
    .A2(_044_),
    .ZN(_047_));
 INV_X4 _357_ (.A(\dpath.a_lt_b$in1[2] ),
    .ZN(_048_));
 NAND2_X4 _358_ (.A1(_048_),
    .A2(\dpath.a_lt_b$in0[2] ),
    .ZN(_049_));
 INV_X2 _359_ (.A(\dpath.a_lt_b$in0[2] ),
    .ZN(_050_));
 NAND2_X4 _360_ (.A1(_050_),
    .A2(\dpath.a_lt_b$in1[2] ),
    .ZN(_051_));
 NAND2_X4 _361_ (.A1(_049_),
    .A2(_051_),
    .ZN(_052_));
 NOR2_X4 _362_ (.A1(_052_),
    .A2(_047_),
    .ZN(_053_));
 NAND2_X4 _363_ (.A1(_042_),
    .A2(_053_),
    .ZN(_054_));
 INV_X2 _364_ (.A(_046_),
    .ZN(_055_));
 OAI21_X1 _365_ (.A(_044_),
    .B1(_055_),
    .B2(_049_),
    .ZN(_056_));
 INV_X2 _366_ (.A(_056_),
    .ZN(_057_));
 NAND2_X4 _367_ (.A1(_054_),
    .A2(_057_),
    .ZN(_058_));
 BUF_X8 _368_ (.A(\dpath.a_lt_b$in0[5] ),
    .Z(_059_));
 XNOR2_X2 _369_ (.A(_059_),
    .B(\dpath.a_lt_b$in1[5] ),
    .ZN(_060_));
 XNOR2_X2 _370_ (.A(\dpath.a_lt_b$in1[4] ),
    .B(\dpath.a_lt_b$in0[4] ),
    .ZN(_061_));
 NAND2_X2 _371_ (.A1(_061_),
    .A2(_060_),
    .ZN(_062_));
 XNOR2_X2 _372_ (.A(\dpath.a_lt_b$in0[7] ),
    .B(\dpath.a_lt_b$in1[7] ),
    .ZN(_063_));
 XNOR2_X2 _373_ (.A(\dpath.a_lt_b$in0[6] ),
    .B(\dpath.a_lt_b$in1[6] ),
    .ZN(_064_));
 NAND2_X4 _374_ (.A1(_064_),
    .A2(_063_),
    .ZN(_065_));
 NOR2_X4 _375_ (.A1(_065_),
    .A2(_062_),
    .ZN(_066_));
 NAND2_X4 _376_ (.A1(_066_),
    .A2(_058_),
    .ZN(_067_));
 INV_X2 _377_ (.A(\dpath.a_lt_b$in1[4] ),
    .ZN(_068_));
 NAND2_X1 _378_ (.A1(_068_),
    .A2(\dpath.a_lt_b$in0[4] ),
    .ZN(_069_));
 INV_X2 _379_ (.A(_059_),
    .ZN(_070_));
 OAI21_X4 _380_ (.A(_069_),
    .B1(\dpath.a_lt_b$in1[5] ),
    .B2(_070_),
    .ZN(_071_));
 INV_X2 _381_ (.A(\dpath.a_lt_b$in1[5] ),
    .ZN(_072_));
 NOR2_X4 _382_ (.A1(_072_),
    .A2(_059_),
    .ZN(_073_));
 INV_X2 _383_ (.A(_073_),
    .ZN(_074_));
 NAND2_X2 _384_ (.A1(_071_),
    .A2(_074_),
    .ZN(_075_));
 NOR2_X4 _385_ (.A1(_075_),
    .A2(_065_),
    .ZN(_076_));
 INV_X2 _386_ (.A(\dpath.a_lt_b$in1[7] ),
    .ZN(_077_));
 NAND2_X1 _387_ (.A1(_077_),
    .A2(\dpath.a_lt_b$in0[7] ),
    .ZN(_078_));
 INV_X4 _388_ (.A(_063_),
    .ZN(_079_));
 INV_X2 _389_ (.A(\dpath.a_lt_b$in1[6] ),
    .ZN(_080_));
 NAND2_X1 _390_ (.A1(_080_),
    .A2(\dpath.a_lt_b$in0[6] ),
    .ZN(_081_));
 OAI21_X2 _391_ (.A(_078_),
    .B1(_079_),
    .B2(_081_),
    .ZN(_082_));
 NOR2_X4 _392_ (.A1(_076_),
    .A2(_082_),
    .ZN(_083_));
 NAND2_X4 _393_ (.A1(_067_),
    .A2(_083_),
    .ZN(_084_));
 INV_X4 _394_ (.A(\dpath.a_lt_b$in1[11] ),
    .ZN(_085_));
 XNOR2_X2 _395_ (.A(_085_),
    .B(\dpath.a_lt_b$in0[11] ),
    .ZN(_086_));
 INV_X4 _396_ (.A(\dpath.a_lt_b$in1[10] ),
    .ZN(_087_));
 XNOR2_X2 _397_ (.A(_087_),
    .B(\dpath.a_lt_b$in0[10] ),
    .ZN(_088_));
 NOR2_X4 _398_ (.A1(_086_),
    .A2(_088_),
    .ZN(_089_));
 XNOR2_X2 _399_ (.A(\dpath.a_lt_b$in0[9] ),
    .B(\dpath.a_lt_b$in1[9] ),
    .ZN(_090_));
 XNOR2_X2 _400_ (.A(\dpath.a_lt_b$in1[8] ),
    .B(\dpath.a_lt_b$in0[8] ),
    .ZN(_091_));
 NAND2_X1 _401_ (.A1(_090_),
    .A2(_091_),
    .ZN(_092_));
 INV_X2 _402_ (.A(_092_),
    .ZN(_093_));
 AND2_X2 _403_ (.A1(_089_),
    .A2(_093_),
    .ZN(_094_));
 NAND2_X4 _404_ (.A1(_084_),
    .A2(_094_),
    .ZN(_095_));
 NAND2_X1 _405_ (.A1(_085_),
    .A2(\dpath.a_lt_b$in0[11] ),
    .ZN(_096_));
 NAND2_X1 _406_ (.A1(_087_),
    .A2(\dpath.a_lt_b$in0[10] ),
    .ZN(_097_));
 OAI21_X2 _407_ (.A(_096_),
    .B1(_086_),
    .B2(_097_),
    .ZN(_098_));
 INV_X2 _408_ (.A(\dpath.a_lt_b$in0[9] ),
    .ZN(_099_));
 NOR2_X1 _409_ (.A1(_099_),
    .A2(\dpath.a_lt_b$in1[9] ),
    .ZN(_100_));
 INV_X2 _410_ (.A(\dpath.a_lt_b$in1[8] ),
    .ZN(_101_));
 AND2_X2 _411_ (.A1(_101_),
    .A2(\dpath.a_lt_b$in0[8] ),
    .ZN(_102_));
 AOI21_X4 _412_ (.A(_100_),
    .B1(_090_),
    .B2(_102_),
    .ZN(_103_));
 INV_X2 _413_ (.A(_103_),
    .ZN(_104_));
 AOI21_X4 _414_ (.A(_098_),
    .B1(_104_),
    .B2(_089_),
    .ZN(_105_));
 NAND2_X4 _415_ (.A1(_095_),
    .A2(_105_),
    .ZN(_106_));
 XNOR2_X2 _416_ (.A(\dpath.a_lt_b$in1[12] ),
    .B(\dpath.a_lt_b$in0[12] ),
    .ZN(_107_));
 INV_X2 _417_ (.A(_107_),
    .ZN(_108_));
 INV_X4 _418_ (.A(\dpath.a_lt_b$in1[13] ),
    .ZN(_109_));
 XNOR2_X2 _419_ (.A(_109_),
    .B(\dpath.a_lt_b$in0[13] ),
    .ZN(_110_));
 NOR2_X4 _420_ (.A1(_108_),
    .A2(_110_),
    .ZN(_111_));
 NAND2_X4 _421_ (.A1(_106_),
    .A2(_111_),
    .ZN(_112_));
 NAND2_X1 _422_ (.A1(_109_),
    .A2(\dpath.a_lt_b$in0[13] ),
    .ZN(_113_));
 INV_X1 _423_ (.A(\dpath.a_lt_b$in1[12] ),
    .ZN(_114_));
 NAND2_X1 _424_ (.A1(_114_),
    .A2(\dpath.a_lt_b$in0[12] ),
    .ZN(_115_));
 OAI21_X1 _425_ (.A(_113_),
    .B1(_110_),
    .B2(_115_),
    .ZN(_116_));
 INV_X1 _426_ (.A(_116_),
    .ZN(_117_));
 NAND2_X4 _427_ (.A1(_112_),
    .A2(_117_),
    .ZN(_118_));
 INV_X1 _428_ (.A(\dpath.a_lt_b$in1[14] ),
    .ZN(_119_));
 XNOR2_X1 _429_ (.A(_119_),
    .B(\dpath.a_lt_b$in0[14] ),
    .ZN(_120_));
 INV_X1 _430_ (.A(_120_),
    .ZN(_121_));
 NAND2_X4 _431_ (.A1(_118_),
    .A2(_121_),
    .ZN(_122_));
 NAND2_X1 _432_ (.A1(_119_),
    .A2(\dpath.a_lt_b$in0[14] ),
    .ZN(_123_));
 NAND2_X4 _433_ (.A1(_122_),
    .A2(_123_),
    .ZN(_124_));
 INV_X1 _434_ (.A(\dpath.a_lt_b$in1[15] ),
    .ZN(_125_));
 XNOR2_X2 _435_ (.A(_125_),
    .B(\dpath.a_lt_b$in0[15] ),
    .ZN(_126_));
 INV_X1 _436_ (.A(_126_),
    .ZN(_127_));
 NAND2_X4 _437_ (.A1(_124_),
    .A2(_127_),
    .ZN(_128_));
 NAND3_X2 _438_ (.A1(_122_),
    .A2(_123_),
    .A3(_126_),
    .ZN(_129_));
 AND2_X2 _439_ (.A1(_128_),
    .A2(_129_),
    .ZN(resp_msg[15]));
 XNOR2_X1 _440_ (.A(\dpath.a_lt_b$in1[1] ),
    .B(_037_),
    .ZN(_130_));
 INV_X1 _441_ (.A(_040_),
    .ZN(_131_));
 XNOR2_X1 _442_ (.A(_130_),
    .B(_131_),
    .ZN(_132_));
 INV_X1 _443_ (.A(_132_),
    .ZN(resp_msg[1]));
 INV_X1 _444_ (.A(_052_),
    .ZN(_133_));
 XNOR2_X1 _445_ (.A(_042_),
    .B(_133_),
    .ZN(_134_));
 INV_X1 _446_ (.A(_134_),
    .ZN(resp_msg[2]));
 NAND2_X1 _447_ (.A1(_042_),
    .A2(_133_),
    .ZN(_135_));
 NAND2_X1 _448_ (.A1(_135_),
    .A2(_049_),
    .ZN(_136_));
 XNOR2_X1 _449_ (.A(_136_),
    .B(_047_),
    .ZN(resp_msg[3]));
 XNOR2_X1 _450_ (.A(_058_),
    .B(_061_),
    .ZN(_137_));
 INV_X1 _451_ (.A(_137_),
    .ZN(resp_msg[4]));
 NAND2_X1 _452_ (.A1(_058_),
    .A2(_061_),
    .ZN(_138_));
 NAND2_X1 _453_ (.A1(_138_),
    .A2(_069_),
    .ZN(_139_));
 XOR2_X1 _454_ (.A(_139_),
    .B(_060_),
    .Z(resp_msg[5]));
 INV_X1 _455_ (.A(_071_),
    .ZN(_140_));
 AOI21_X4 _456_ (.A(_073_),
    .B1(_138_),
    .B2(_140_),
    .ZN(_141_));
 XNOR2_X2 _457_ (.A(_141_),
    .B(_064_),
    .ZN(_142_));
 INV_X2 _458_ (.A(_142_),
    .ZN(resp_msg[6]));
 NAND2_X1 _459_ (.A1(_141_),
    .A2(_064_),
    .ZN(_143_));
 NAND2_X1 _460_ (.A1(_143_),
    .A2(_081_),
    .ZN(_144_));
 XNOR2_X2 _461_ (.A(_144_),
    .B(_079_),
    .ZN(resp_msg[7]));
 XNOR2_X1 _462_ (.A(_084_),
    .B(_091_),
    .ZN(_145_));
 INV_X1 _463_ (.A(_145_),
    .ZN(resp_msg[8]));
 AOI21_X1 _464_ (.A(_102_),
    .B1(_084_),
    .B2(_091_),
    .ZN(_146_));
 XNOR2_X2 _465_ (.A(_146_),
    .B(_090_),
    .ZN(resp_msg[9]));
 NAND2_X1 _466_ (.A1(_084_),
    .A2(_093_),
    .ZN(_147_));
 NAND2_X4 _467_ (.A1(_147_),
    .A2(_103_),
    .ZN(_148_));
 INV_X1 _468_ (.A(_088_),
    .ZN(_149_));
 XNOR2_X2 _469_ (.A(_148_),
    .B(_149_),
    .ZN(_150_));
 INV_X2 _470_ (.A(_150_),
    .ZN(resp_msg[10]));
 NAND2_X4 _471_ (.A1(_148_),
    .A2(_149_),
    .ZN(_151_));
 NAND2_X4 _472_ (.A1(_151_),
    .A2(_097_),
    .ZN(_152_));
 XNOR2_X2 _473_ (.A(_152_),
    .B(_086_),
    .ZN(resp_msg[11]));
 XNOR2_X2 _474_ (.A(_106_),
    .B(_107_),
    .ZN(_153_));
 INV_X2 _475_ (.A(_153_),
    .ZN(resp_msg[12]));
 NAND2_X4 _476_ (.A1(_106_),
    .A2(_107_),
    .ZN(_154_));
 NAND2_X4 _477_ (.A1(_154_),
    .A2(_115_),
    .ZN(_155_));
 XNOR2_X2 _478_ (.A(_110_),
    .B(_155_),
    .ZN(resp_msg[13]));
 XNOR2_X2 _479_ (.A(_118_),
    .B(_121_),
    .ZN(_156_));
 INV_X2 _480_ (.A(_156_),
    .ZN(resp_msg[14]));
 XNOR2_X1 _481_ (.A(_039_),
    .B(\dpath.a_lt_b$in0[0] ),
    .ZN(resp_msg[0]));
 NAND4_X1 _482_ (.A1(_119_),
    .A2(_125_),
    .A3(_039_),
    .A4(_036_),
    .ZN(_157_));
 NAND3_X1 _483_ (.A1(_087_),
    .A2(_085_),
    .A3(_114_),
    .ZN(_158_));
 NOR3_X1 _484_ (.A1(_157_),
    .A2(\dpath.a_lt_b$in1[13] ),
    .A3(_158_),
    .ZN(_159_));
 INV_X1 _485_ (.A(\dpath.a_lt_b$in1[9] ),
    .ZN(_160_));
 NAND4_X1 _486_ (.A1(_080_),
    .A2(_077_),
    .A3(_101_),
    .A4(_160_),
    .ZN(_161_));
 NAND4_X1 _487_ (.A1(_048_),
    .A2(_043_),
    .A3(_068_),
    .A4(_072_),
    .ZN(_162_));
 NOR2_X1 _488_ (.A1(_161_),
    .A2(_162_),
    .ZN(_163_));
 NAND2_X1 _489_ (.A1(_159_),
    .A2(_163_),
    .ZN(_164_));
 INV_X1 _490_ (.A(_164_),
    .ZN(_165_));
 BUF_X1 _491_ (.A(\ctrl.state.out[2] ),
    .Z(_166_));
 INV_X1 _492_ (.A(_166_),
    .ZN(_167_));
 OR2_X1 _493_ (.A1(_167_),
    .A2(reset),
    .ZN(_168_));
 CLKBUF_X1 _494_ (.A(req_rdy),
    .Z(_169_));
 BUF_X1 _495_ (.A(_169_),
    .Z(_170_));
 BUF_X1 _496_ (.A(_170_),
    .Z(_171_));
 NAND2_X1 _497_ (.A1(_171_),
    .A2(req_val),
    .ZN(_172_));
 OAI22_X1 _498_ (.A1(_165_),
    .A2(_168_),
    .B1(reset),
    .B2(_172_),
    .ZN(_002_));
 BUF_X1 _499_ (.A(_003_),
    .Z(_173_));
 AND3_X1 _500_ (.A1(_167_),
    .A2(_173_),
    .A3(\ctrl.state.out[1] ),
    .ZN(resp_val));
 AOI21_X1 _501_ (.A(reset),
    .B1(resp_val),
    .B2(resp_rdy),
    .ZN(_174_));
 BUF_X1 _502_ (.A(_170_),
    .Z(_175_));
 INV_X1 _503_ (.A(_175_),
    .ZN(_176_));
 OAI21_X1 _504_ (.A(_174_),
    .B1(_176_),
    .B2(req_val),
    .ZN(_000_));
 NAND2_X1 _505_ (.A1(_174_),
    .A2(\ctrl.state.out[1] ),
    .ZN(_177_));
 OAI21_X1 _506_ (.A(_177_),
    .B1(_164_),
    .B2(_168_),
    .ZN(_001_));
 NAND2_X1 _507_ (.A1(_125_),
    .A2(\dpath.a_lt_b$in0[15] ),
    .ZN(_178_));
 OAI21_X1 _508_ (.A(_178_),
    .B1(_126_),
    .B2(_123_),
    .ZN(_179_));
 NOR2_X4 _509_ (.A1(_120_),
    .A2(_126_),
    .ZN(_180_));
 AOI21_X1 _510_ (.A(_179_),
    .B1(_116_),
    .B2(_180_),
    .ZN(_181_));
 NAND2_X1 _511_ (.A1(_111_),
    .A2(_180_),
    .ZN(_182_));
 OAI21_X1 _512_ (.A(_181_),
    .B1(_105_),
    .B2(_182_),
    .ZN(_183_));
 INV_X4 _513_ (.A(_183_),
    .ZN(_184_));
 INV_X2 _514_ (.A(_182_),
    .ZN(_185_));
 NAND3_X4 _515_ (.A1(_084_),
    .A2(_094_),
    .A3(_185_),
    .ZN(_186_));
 NAND3_X2 _516_ (.A1(_184_),
    .A2(_186_),
    .A3(_166_),
    .ZN(_187_));
 NAND2_X4 _517_ (.A1(_187_),
    .A2(_173_),
    .ZN(_188_));
 BUF_X2 _518_ (.A(_188_),
    .Z(_189_));
 MUX2_X1 _519_ (.A(\dpath.a_lt_b$in0[0] ),
    .B(req_msg[0]),
    .S(_170_),
    .Z(_190_));
 NAND2_X1 _520_ (.A1(_189_),
    .A2(_190_),
    .ZN(_191_));
 BUF_X2 _521_ (.A(_188_),
    .Z(_192_));
 OAI21_X1 _522_ (.A(_191_),
    .B1(_039_),
    .B2(_192_),
    .ZN(_004_));
 MUX2_X1 _523_ (.A(_037_),
    .B(req_msg[1]),
    .S(_170_),
    .Z(_193_));
 NAND2_X1 _524_ (.A1(_189_),
    .A2(_193_),
    .ZN(_194_));
 OAI21_X1 _525_ (.A(_194_),
    .B1(_036_),
    .B2(_192_),
    .ZN(_005_));
 NAND2_X1 _526_ (.A1(_170_),
    .A2(req_msg[2]),
    .ZN(_195_));
 OAI21_X1 _527_ (.A(_195_),
    .B1(_171_),
    .B2(_050_),
    .ZN(_196_));
 NAND2_X1 _528_ (.A1(_189_),
    .A2(_196_),
    .ZN(_197_));
 OAI21_X1 _529_ (.A(_197_),
    .B1(_048_),
    .B2(_192_),
    .ZN(_006_));
 NAND2_X1 _530_ (.A1(_170_),
    .A2(req_msg[3]),
    .ZN(_198_));
 OAI21_X1 _531_ (.A(_198_),
    .B1(_171_),
    .B2(_045_),
    .ZN(_199_));
 NAND2_X1 _532_ (.A1(_189_),
    .A2(_199_),
    .ZN(_200_));
 OAI21_X1 _533_ (.A(_200_),
    .B1(_043_),
    .B2(_192_),
    .ZN(_007_));
 BUF_X2 _534_ (.A(_188_),
    .Z(_201_));
 BUF_X1 _535_ (.A(_169_),
    .Z(_202_));
 MUX2_X1 _536_ (.A(\dpath.a_lt_b$in0[4] ),
    .B(req_msg[4]),
    .S(_202_),
    .Z(_203_));
 NAND2_X1 _537_ (.A1(_201_),
    .A2(_203_),
    .ZN(_204_));
 OAI21_X1 _538_ (.A(_204_),
    .B1(_068_),
    .B2(_192_),
    .ZN(_008_));
 NAND2_X1 _539_ (.A1(_170_),
    .A2(req_msg[5]),
    .ZN(_205_));
 OAI21_X1 _540_ (.A(_205_),
    .B1(_170_),
    .B2(_070_),
    .ZN(_206_));
 NAND2_X1 _541_ (.A1(_201_),
    .A2(_206_),
    .ZN(_207_));
 OAI21_X1 _542_ (.A(_207_),
    .B1(_072_),
    .B2(_192_),
    .ZN(_009_));
 MUX2_X1 _543_ (.A(\dpath.a_lt_b$in0[6] ),
    .B(req_msg[6]),
    .S(_202_),
    .Z(_208_));
 NAND2_X1 _544_ (.A1(_201_),
    .A2(_208_),
    .ZN(_209_));
 OAI21_X1 _545_ (.A(_209_),
    .B1(_080_),
    .B2(_192_),
    .ZN(_010_));
 MUX2_X1 _546_ (.A(\dpath.a_lt_b$in0[7] ),
    .B(req_msg[7]),
    .S(_202_),
    .Z(_210_));
 NAND2_X1 _547_ (.A1(_201_),
    .A2(_210_),
    .ZN(_211_));
 OAI21_X1 _548_ (.A(_211_),
    .B1(_077_),
    .B2(_192_),
    .ZN(_011_));
 MUX2_X1 _549_ (.A(\dpath.a_lt_b$in0[8] ),
    .B(req_msg[8]),
    .S(_202_),
    .Z(_212_));
 NAND2_X1 _550_ (.A1(_201_),
    .A2(_212_),
    .ZN(_213_));
 OAI21_X1 _551_ (.A(_213_),
    .B1(_101_),
    .B2(_192_),
    .ZN(_012_));
 NAND2_X1 _552_ (.A1(_170_),
    .A2(req_msg[9]),
    .ZN(_214_));
 OAI21_X1 _553_ (.A(_214_),
    .B1(_170_),
    .B2(_099_),
    .ZN(_215_));
 NAND2_X1 _554_ (.A1(_201_),
    .A2(_215_),
    .ZN(_216_));
 OAI21_X1 _555_ (.A(_216_),
    .B1(_160_),
    .B2(_192_),
    .ZN(_013_));
 MUX2_X1 _556_ (.A(\dpath.a_lt_b$in0[10] ),
    .B(req_msg[10]),
    .S(_202_),
    .Z(_217_));
 NAND2_X1 _557_ (.A1(_201_),
    .A2(_217_),
    .ZN(_218_));
 OAI21_X1 _558_ (.A(_218_),
    .B1(_087_),
    .B2(_189_),
    .ZN(_014_));
 MUX2_X1 _559_ (.A(\dpath.a_lt_b$in0[11] ),
    .B(req_msg[11]),
    .S(_202_),
    .Z(_219_));
 NAND2_X1 _560_ (.A1(_201_),
    .A2(_219_),
    .ZN(_220_));
 OAI21_X1 _561_ (.A(_220_),
    .B1(_085_),
    .B2(_189_),
    .ZN(_015_));
 MUX2_X1 _562_ (.A(\dpath.a_lt_b$in0[12] ),
    .B(req_msg[12]),
    .S(_202_),
    .Z(_221_));
 NAND2_X1 _563_ (.A1(_201_),
    .A2(_221_),
    .ZN(_222_));
 OAI21_X1 _564_ (.A(_222_),
    .B1(_114_),
    .B2(_189_),
    .ZN(_016_));
 MUX2_X1 _565_ (.A(\dpath.a_lt_b$in0[13] ),
    .B(req_msg[13]),
    .S(_202_),
    .Z(_223_));
 NAND2_X1 _566_ (.A1(_201_),
    .A2(_223_),
    .ZN(_224_));
 OAI21_X1 _567_ (.A(_224_),
    .B1(_109_),
    .B2(_189_),
    .ZN(_017_));
 MUX2_X1 _568_ (.A(\dpath.a_lt_b$in0[14] ),
    .B(req_msg[14]),
    .S(_202_),
    .Z(_225_));
 NAND2_X1 _569_ (.A1(_188_),
    .A2(_225_),
    .ZN(_226_));
 OAI21_X1 _570_ (.A(_226_),
    .B1(_119_),
    .B2(_189_),
    .ZN(_018_));
 MUX2_X1 _571_ (.A(\dpath.a_lt_b$in0[15] ),
    .B(req_msg[15]),
    .S(_202_),
    .Z(_227_));
 NAND2_X1 _572_ (.A1(_188_),
    .A2(_227_),
    .ZN(_228_));
 OAI21_X1 _573_ (.A(_228_),
    .B1(_125_),
    .B2(_189_),
    .ZN(_019_));
 NAND2_X4 _574_ (.A1(_184_),
    .A2(_186_),
    .ZN(_229_));
 NAND3_X4 _575_ (.A1(_229_),
    .A2(_166_),
    .A3(_173_),
    .ZN(_230_));
 INV_X8 _576_ (.A(_230_),
    .ZN(_231_));
 NAND2_X1 _577_ (.A1(_231_),
    .A2(resp_msg[0]),
    .ZN(_232_));
 NAND4_X4 _578_ (.A1(_184_),
    .A2(_186_),
    .A3(_166_),
    .A4(_173_),
    .ZN(_233_));
 BUF_X8 _579_ (.A(_233_),
    .Z(_234_));
 OAI21_X1 _580_ (.A(_232_),
    .B1(_234_),
    .B2(_039_),
    .ZN(_235_));
 NOR2_X1 _581_ (.A1(_167_),
    .A2(_169_),
    .ZN(_236_));
 BUF_X1 _582_ (.A(_236_),
    .Z(_237_));
 NAND2_X1 _583_ (.A1(_235_),
    .A2(_237_),
    .ZN(_238_));
 NAND2_X1 _584_ (.A1(_175_),
    .A2(req_msg[16]),
    .ZN(_239_));
 NOR2_X1 _585_ (.A1(_166_),
    .A2(_169_),
    .ZN(_240_));
 BUF_X1 _586_ (.A(_240_),
    .Z(_241_));
 NAND2_X1 _587_ (.A1(_241_),
    .A2(\dpath.a_lt_b$in0[0] ),
    .ZN(_242_));
 NAND3_X1 _588_ (.A1(_238_),
    .A2(_239_),
    .A3(_242_),
    .ZN(_020_));
 OAI22_X1 _589_ (.A1(_234_),
    .A2(_036_),
    .B1(_230_),
    .B2(_132_),
    .ZN(_243_));
 NAND2_X1 _590_ (.A1(_243_),
    .A2(_237_),
    .ZN(_244_));
 NAND2_X1 _591_ (.A1(_175_),
    .A2(req_msg[17]),
    .ZN(_245_));
 NAND2_X1 _592_ (.A1(_241_),
    .A2(_037_),
    .ZN(_246_));
 NAND3_X1 _593_ (.A1(_244_),
    .A2(_245_),
    .A3(_246_),
    .ZN(_021_));
 OAI22_X1 _594_ (.A1(_234_),
    .A2(_048_),
    .B1(_230_),
    .B2(_134_),
    .ZN(_247_));
 NAND2_X1 _595_ (.A1(_247_),
    .A2(_237_),
    .ZN(_248_));
 NAND2_X1 _596_ (.A1(req_msg[18]),
    .A2(_175_),
    .ZN(_249_));
 NAND2_X1 _597_ (.A1(_241_),
    .A2(\dpath.a_lt_b$in0[2] ),
    .ZN(_250_));
 NAND3_X2 _598_ (.A1(_248_),
    .A2(_249_),
    .A3(_250_),
    .ZN(_022_));
 NAND2_X1 _599_ (.A1(_231_),
    .A2(resp_msg[3]),
    .ZN(_251_));
 OAI21_X1 _600_ (.A(_251_),
    .B1(_234_),
    .B2(_043_),
    .ZN(_252_));
 NAND2_X1 _601_ (.A1(_252_),
    .A2(_237_),
    .ZN(_253_));
 NAND2_X1 _602_ (.A1(req_msg[19]),
    .A2(_175_),
    .ZN(_254_));
 NAND2_X1 _603_ (.A1(_241_),
    .A2(\dpath.a_lt_b$in0[3] ),
    .ZN(_255_));
 NAND3_X1 _604_ (.A1(_253_),
    .A2(_254_),
    .A3(_255_),
    .ZN(_023_));
 OAI22_X1 _605_ (.A1(_234_),
    .A2(_068_),
    .B1(_230_),
    .B2(_137_),
    .ZN(_256_));
 NAND2_X1 _606_ (.A1(_256_),
    .A2(_237_),
    .ZN(_257_));
 NAND2_X1 _607_ (.A1(req_msg[20]),
    .A2(_175_),
    .ZN(_258_));
 NAND2_X1 _608_ (.A1(_241_),
    .A2(\dpath.a_lt_b$in0[4] ),
    .ZN(_259_));
 NAND3_X1 _609_ (.A1(_257_),
    .A2(_258_),
    .A3(_259_),
    .ZN(_024_));
 NAND2_X1 _610_ (.A1(_231_),
    .A2(resp_msg[5]),
    .ZN(_260_));
 OAI21_X1 _611_ (.A(_260_),
    .B1(_234_),
    .B2(_072_),
    .ZN(_261_));
 NAND2_X1 _612_ (.A1(_261_),
    .A2(_237_),
    .ZN(_262_));
 NAND2_X1 _613_ (.A1(req_msg[21]),
    .A2(_175_),
    .ZN(_263_));
 NAND2_X1 _614_ (.A1(_241_),
    .A2(_059_),
    .ZN(_264_));
 NAND3_X1 _615_ (.A1(_262_),
    .A2(_263_),
    .A3(_264_),
    .ZN(_025_));
 OAI22_X1 _616_ (.A1(_234_),
    .A2(_080_),
    .B1(_230_),
    .B2(_142_),
    .ZN(_265_));
 NAND2_X1 _617_ (.A1(_265_),
    .A2(_236_),
    .ZN(_266_));
 NAND2_X1 _618_ (.A1(req_msg[22]),
    .A2(_175_),
    .ZN(_267_));
 NAND2_X1 _619_ (.A1(_241_),
    .A2(\dpath.a_lt_b$in0[6] ),
    .ZN(_268_));
 NAND3_X1 _620_ (.A1(_266_),
    .A2(_267_),
    .A3(_268_),
    .ZN(_026_));
 NAND2_X1 _621_ (.A1(resp_msg[7]),
    .A2(_231_),
    .ZN(_269_));
 OAI21_X1 _622_ (.A(_269_),
    .B1(_077_),
    .B2(_233_),
    .ZN(_270_));
 NAND2_X1 _623_ (.A1(_270_),
    .A2(_236_),
    .ZN(_271_));
 NAND2_X1 _624_ (.A1(req_msg[23]),
    .A2(_175_),
    .ZN(_272_));
 NAND2_X1 _625_ (.A1(_241_),
    .A2(\dpath.a_lt_b$in0[7] ),
    .ZN(_273_));
 NAND3_X1 _626_ (.A1(_271_),
    .A2(_272_),
    .A3(_273_),
    .ZN(_027_));
 OAI22_X1 _627_ (.A1(_233_),
    .A2(_101_),
    .B1(_230_),
    .B2(_145_),
    .ZN(_274_));
 NAND2_X1 _628_ (.A1(_274_),
    .A2(_236_),
    .ZN(_275_));
 NAND2_X1 _629_ (.A1(req_msg[24]),
    .A2(_175_),
    .ZN(_276_));
 NAND2_X1 _630_ (.A1(_241_),
    .A2(\dpath.a_lt_b$in0[8] ),
    .ZN(_277_));
 NAND3_X1 _631_ (.A1(_275_),
    .A2(_276_),
    .A3(_277_),
    .ZN(_028_));
 NAND2_X1 _632_ (.A1(_231_),
    .A2(resp_msg[9]),
    .ZN(_278_));
 OAI21_X1 _633_ (.A(_278_),
    .B1(_234_),
    .B2(_160_),
    .ZN(_279_));
 NAND2_X1 _634_ (.A1(_279_),
    .A2(_236_),
    .ZN(_280_));
 NAND2_X1 _635_ (.A1(req_msg[25]),
    .A2(_171_),
    .ZN(_281_));
 NAND2_X1 _636_ (.A1(_241_),
    .A2(\dpath.a_lt_b$in0[9] ),
    .ZN(_282_));
 NAND3_X1 _637_ (.A1(_280_),
    .A2(_281_),
    .A3(_282_),
    .ZN(_029_));
 OAI22_X1 _638_ (.A1(_150_),
    .A2(_230_),
    .B1(_233_),
    .B2(_087_),
    .ZN(_283_));
 NAND2_X1 _639_ (.A1(_283_),
    .A2(_236_),
    .ZN(_284_));
 NAND2_X1 _640_ (.A1(req_msg[26]),
    .A2(_171_),
    .ZN(_285_));
 NAND2_X1 _641_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[10] ),
    .ZN(_286_));
 NAND3_X1 _642_ (.A1(_284_),
    .A2(_285_),
    .A3(_286_),
    .ZN(_030_));
 NAND2_X1 _643_ (.A1(resp_msg[11]),
    .A2(_231_),
    .ZN(_287_));
 OAI21_X1 _644_ (.A(_287_),
    .B1(_085_),
    .B2(_234_),
    .ZN(_288_));
 NAND2_X1 _645_ (.A1(_288_),
    .A2(_237_),
    .ZN(_289_));
 AND2_X1 _646_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[11] ),
    .ZN(_290_));
 AOI21_X1 _647_ (.A(_290_),
    .B1(req_msg[27]),
    .B2(_171_),
    .ZN(_291_));
 NAND2_X1 _648_ (.A1(_289_),
    .A2(_291_),
    .ZN(_031_));
 OAI22_X1 _649_ (.A1(_153_),
    .A2(_230_),
    .B1(_233_),
    .B2(_114_),
    .ZN(_292_));
 NAND2_X1 _650_ (.A1(_292_),
    .A2(_236_),
    .ZN(_293_));
 NAND2_X1 _651_ (.A1(req_msg[28]),
    .A2(_171_),
    .ZN(_294_));
 NAND2_X1 _652_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[12] ),
    .ZN(_295_));
 NAND3_X1 _653_ (.A1(_293_),
    .A2(_294_),
    .A3(_295_),
    .ZN(_032_));
 NAND2_X1 _654_ (.A1(resp_msg[13]),
    .A2(_231_),
    .ZN(_296_));
 OAI21_X1 _655_ (.A(_296_),
    .B1(_109_),
    .B2(_234_),
    .ZN(_297_));
 NAND2_X1 _656_ (.A1(_297_),
    .A2(_237_),
    .ZN(_298_));
 AND2_X1 _657_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[13] ),
    .ZN(_299_));
 AOI21_X1 _658_ (.A(_299_),
    .B1(req_msg[29]),
    .B2(_171_),
    .ZN(_300_));
 NAND2_X1 _659_ (.A1(_298_),
    .A2(_300_),
    .ZN(_033_));
 OAI22_X1 _660_ (.A1(_156_),
    .A2(_230_),
    .B1(_233_),
    .B2(_119_),
    .ZN(_301_));
 NAND2_X1 _661_ (.A1(_301_),
    .A2(_237_),
    .ZN(_302_));
 AND2_X1 _662_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[14] ),
    .ZN(_303_));
 AOI21_X1 _663_ (.A(_303_),
    .B1(req_msg[30]),
    .B2(_171_),
    .ZN(_304_));
 NAND2_X1 _664_ (.A1(_302_),
    .A2(_304_),
    .ZN(_034_));
 NAND3_X1 _665_ (.A1(_128_),
    .A2(_129_),
    .A3(_231_),
    .ZN(_305_));
 OR2_X2 _666_ (.A1(_233_),
    .A2(_125_),
    .ZN(_306_));
 NAND2_X1 _667_ (.A1(_305_),
    .A2(_306_),
    .ZN(_307_));
 NAND2_X1 _668_ (.A1(_307_),
    .A2(_237_),
    .ZN(_308_));
 AND2_X1 _669_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[15] ),
    .ZN(_309_));
 AOI21_X1 _670_ (.A(_309_),
    .B1(req_msg[31]),
    .B2(_171_),
    .ZN(_310_));
 NAND2_X1 _671_ (.A1(_308_),
    .A2(_310_),
    .ZN(_035_));
 DFF_X1 _672_ (.D(_000_),
    .CK(clknet_2_2__leaf_clk),
    .Q(req_rdy),
    .QN(_003_));
 DFF_X1 _673_ (.D(_001_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\ctrl.state.out[1] ),
    .QN(_311_));
 DFF_X1 _674_ (.D(_002_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\ctrl.state.out[2] ),
    .QN(_312_));
 DFF_X1 _675_ (.D(_004_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in1[0] ),
    .QN(_313_));
 DFF_X1 _676_ (.D(_005_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in1[1] ),
    .QN(_314_));
 DFF_X1 _677_ (.D(_006_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in1[2] ),
    .QN(_315_));
 DFF_X1 _678_ (.D(_007_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in1[3] ),
    .QN(_316_));
 DFF_X1 _679_ (.D(_008_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in1[4] ),
    .QN(_317_));
 DFF_X1 _680_ (.D(_009_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in1[5] ),
    .QN(_318_));
 DFF_X1 _681_ (.D(_010_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in1[6] ),
    .QN(_319_));
 DFF_X1 _682_ (.D(_011_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in1[7] ),
    .QN(_320_));
 DFF_X1 _683_ (.D(_012_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in1[8] ),
    .QN(_321_));
 DFF_X1 _684_ (.D(_013_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in1[9] ),
    .QN(_322_));
 DFF_X1 _685_ (.D(_014_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in1[10] ),
    .QN(_323_));
 DFF_X1 _686_ (.D(_015_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in1[11] ),
    .QN(_324_));
 DFF_X1 _687_ (.D(_016_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in1[12] ),
    .QN(_325_));
 DFF_X1 _688_ (.D(_017_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in1[13] ),
    .QN(_326_));
 DFF_X1 _689_ (.D(_018_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in1[14] ),
    .QN(_327_));
 DFF_X1 _690_ (.D(_019_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in1[15] ),
    .QN(_328_));
 DFF_X1 _691_ (.D(_020_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in0[0] ),
    .QN(_329_));
 DFF_X1 _692_ (.D(_021_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in0[1] ),
    .QN(_330_));
 DFF_X1 _693_ (.D(_022_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in0[2] ),
    .QN(_331_));
 DFF_X1 _694_ (.D(_023_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in0[3] ),
    .QN(_332_));
 DFF_X1 _695_ (.D(_024_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in0[4] ),
    .QN(_333_));
 DFF_X1 _696_ (.D(_025_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in0[5] ),
    .QN(_334_));
 DFF_X1 _697_ (.D(_026_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in0[6] ),
    .QN(_335_));
 DFF_X1 _698_ (.D(_027_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in0[7] ),
    .QN(_336_));
 DFF_X1 _699_ (.D(_028_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in0[8] ),
    .QN(_337_));
 DFF_X1 _700_ (.D(_029_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in0[9] ),
    .QN(_338_));
 DFF_X1 _701_ (.D(_030_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in0[10] ),
    .QN(_339_));
 DFF_X1 _702_ (.D(_031_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in0[11] ),
    .QN(_340_));
 DFF_X1 _703_ (.D(_032_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in0[12] ),
    .QN(_341_));
 DFF_X1 _704_ (.D(_033_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in0[13] ),
    .QN(_342_));
 DFF_X1 _705_ (.D(_034_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in0[14] ),
    .QN(_343_));
 DFF_X1 _706_ (.D(_035_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in0[15] ),
    .QN(_344_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_113 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_114 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_115 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_116 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_117 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_118 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_119 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_120 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_121 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_122 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_123 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_124 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_125 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_126 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_127 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_128 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_129 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_130 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_131 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_132 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_133 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_134 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_135 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_136 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_137 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_138 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_139 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_140 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_141 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_142 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_143 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_144 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_145 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_146 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_147 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_148 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_149 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_150 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_151 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_152 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_153 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_154 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_155 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_156 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_157 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_158 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_159 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_160 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_161 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_162 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_163 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_164 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_165 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_166 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_167 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_168 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_169 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_170 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_171 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_172 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_173 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_174 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_175 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_176 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_177 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_178 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_179 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_180 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_181 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_182 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_183 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_184 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_185 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_186 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_187 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_188 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_189 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_190 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_191 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_192 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_193 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_194 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_195 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_196 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_197 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_198 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_199 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_200 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_201 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_202 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_203 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_204 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_205 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_206 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_207 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_208 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_209 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_210 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_211 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_212 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_213 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_214 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_215 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_216 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_217 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_218 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_41_219 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_41_220 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_221 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_222 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_223 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_43_224 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_43_225 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_226 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_227 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_228 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_45_229 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_45_230 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_231 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_232 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_233 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_47_234 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_47_235 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_236 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_237 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_238 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_49_239 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_49_240 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_241 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_242 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_243 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_244 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_245 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_246 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_247 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_248 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_53_249 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_53_250 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_251 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_252 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_253 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_55_254 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_55_255 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_256 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_257 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_258 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_259 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_260 ();
 BUF_X4 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 BUF_X4 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 BUF_X4 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 BUF_X4 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 BUF_X4 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 INV_X1 clkload0 (.A(clknet_2_1__leaf_clk));
 INV_X2 clkload1 (.A(clknet_2_3__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X8 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_74 ();
 FILLCELL_X32 FILLER_0_106 ();
 FILLCELL_X8 FILLER_0_138 ();
 FILLCELL_X32 FILLER_0_147 ();
 FILLCELL_X32 FILLER_0_179 ();
 FILLCELL_X8 FILLER_0_211 ();
 FILLCELL_X32 FILLER_0_220 ();
 FILLCELL_X32 FILLER_0_252 ();
 FILLCELL_X8 FILLER_0_284 ();
 FILLCELL_X32 FILLER_0_293 ();
 FILLCELL_X32 FILLER_0_325 ();
 FILLCELL_X8 FILLER_0_357 ();
 FILLCELL_X32 FILLER_0_366 ();
 FILLCELL_X16 FILLER_0_398 ();
 FILLCELL_X4 FILLER_0_414 ();
 FILLCELL_X2 FILLER_0_418 ();
 FILLCELL_X1 FILLER_0_420 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X16 FILLER_1_129 ();
 FILLCELL_X2 FILLER_1_145 ();
 FILLCELL_X32 FILLER_1_148 ();
 FILLCELL_X32 FILLER_1_180 ();
 FILLCELL_X32 FILLER_1_212 ();
 FILLCELL_X32 FILLER_1_244 ();
 FILLCELL_X16 FILLER_1_276 ();
 FILLCELL_X2 FILLER_1_292 ();
 FILLCELL_X32 FILLER_1_295 ();
 FILLCELL_X32 FILLER_1_327 ();
 FILLCELL_X32 FILLER_1_359 ();
 FILLCELL_X16 FILLER_1_391 ();
 FILLCELL_X8 FILLER_1_407 ();
 FILLCELL_X4 FILLER_1_415 ();
 FILLCELL_X2 FILLER_1_419 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X8 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_74 ();
 FILLCELL_X32 FILLER_2_106 ();
 FILLCELL_X32 FILLER_2_138 ();
 FILLCELL_X32 FILLER_2_170 ();
 FILLCELL_X16 FILLER_2_202 ();
 FILLCELL_X2 FILLER_2_218 ();
 FILLCELL_X32 FILLER_2_221 ();
 FILLCELL_X32 FILLER_2_253 ();
 FILLCELL_X32 FILLER_2_285 ();
 FILLCELL_X32 FILLER_2_317 ();
 FILLCELL_X16 FILLER_2_349 ();
 FILLCELL_X2 FILLER_2_365 ();
 FILLCELL_X32 FILLER_2_368 ();
 FILLCELL_X16 FILLER_2_400 ();
 FILLCELL_X4 FILLER_2_416 ();
 FILLCELL_X1 FILLER_2_420 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X16 FILLER_3_129 ();
 FILLCELL_X2 FILLER_3_145 ();
 FILLCELL_X32 FILLER_3_148 ();
 FILLCELL_X32 FILLER_3_180 ();
 FILLCELL_X32 FILLER_3_212 ();
 FILLCELL_X32 FILLER_3_244 ();
 FILLCELL_X16 FILLER_3_276 ();
 FILLCELL_X2 FILLER_3_292 ();
 FILLCELL_X32 FILLER_3_295 ();
 FILLCELL_X32 FILLER_3_327 ();
 FILLCELL_X32 FILLER_3_359 ();
 FILLCELL_X16 FILLER_3_391 ();
 FILLCELL_X8 FILLER_3_407 ();
 FILLCELL_X4 FILLER_3_415 ();
 FILLCELL_X2 FILLER_3_419 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X8 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_74 ();
 FILLCELL_X32 FILLER_4_106 ();
 FILLCELL_X32 FILLER_4_138 ();
 FILLCELL_X32 FILLER_4_170 ();
 FILLCELL_X16 FILLER_4_202 ();
 FILLCELL_X2 FILLER_4_218 ();
 FILLCELL_X32 FILLER_4_221 ();
 FILLCELL_X32 FILLER_4_253 ();
 FILLCELL_X32 FILLER_4_285 ();
 FILLCELL_X32 FILLER_4_317 ();
 FILLCELL_X16 FILLER_4_349 ();
 FILLCELL_X2 FILLER_4_365 ();
 FILLCELL_X32 FILLER_4_368 ();
 FILLCELL_X16 FILLER_4_400 ();
 FILLCELL_X4 FILLER_4_416 ();
 FILLCELL_X1 FILLER_4_420 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X16 FILLER_5_129 ();
 FILLCELL_X2 FILLER_5_145 ();
 FILLCELL_X32 FILLER_5_148 ();
 FILLCELL_X32 FILLER_5_180 ();
 FILLCELL_X32 FILLER_5_212 ();
 FILLCELL_X32 FILLER_5_244 ();
 FILLCELL_X16 FILLER_5_276 ();
 FILLCELL_X2 FILLER_5_292 ();
 FILLCELL_X32 FILLER_5_295 ();
 FILLCELL_X32 FILLER_5_327 ();
 FILLCELL_X32 FILLER_5_359 ();
 FILLCELL_X16 FILLER_5_391 ();
 FILLCELL_X8 FILLER_5_407 ();
 FILLCELL_X4 FILLER_5_415 ();
 FILLCELL_X2 FILLER_5_419 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X8 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_74 ();
 FILLCELL_X32 FILLER_6_106 ();
 FILLCELL_X32 FILLER_6_138 ();
 FILLCELL_X32 FILLER_6_170 ();
 FILLCELL_X16 FILLER_6_202 ();
 FILLCELL_X2 FILLER_6_218 ();
 FILLCELL_X32 FILLER_6_221 ();
 FILLCELL_X32 FILLER_6_253 ();
 FILLCELL_X32 FILLER_6_285 ();
 FILLCELL_X32 FILLER_6_317 ();
 FILLCELL_X16 FILLER_6_349 ();
 FILLCELL_X2 FILLER_6_365 ();
 FILLCELL_X32 FILLER_6_368 ();
 FILLCELL_X16 FILLER_6_400 ();
 FILLCELL_X4 FILLER_6_416 ();
 FILLCELL_X1 FILLER_6_420 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X16 FILLER_7_129 ();
 FILLCELL_X2 FILLER_7_145 ();
 FILLCELL_X32 FILLER_7_148 ();
 FILLCELL_X32 FILLER_7_180 ();
 FILLCELL_X32 FILLER_7_212 ();
 FILLCELL_X32 FILLER_7_244 ();
 FILLCELL_X16 FILLER_7_276 ();
 FILLCELL_X2 FILLER_7_292 ();
 FILLCELL_X32 FILLER_7_295 ();
 FILLCELL_X32 FILLER_7_327 ();
 FILLCELL_X32 FILLER_7_359 ();
 FILLCELL_X16 FILLER_7_391 ();
 FILLCELL_X8 FILLER_7_407 ();
 FILLCELL_X4 FILLER_7_415 ();
 FILLCELL_X2 FILLER_7_419 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X8 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_74 ();
 FILLCELL_X32 FILLER_8_106 ();
 FILLCELL_X32 FILLER_8_138 ();
 FILLCELL_X32 FILLER_8_170 ();
 FILLCELL_X16 FILLER_8_202 ();
 FILLCELL_X2 FILLER_8_218 ();
 FILLCELL_X32 FILLER_8_221 ();
 FILLCELL_X32 FILLER_8_253 ();
 FILLCELL_X32 FILLER_8_285 ();
 FILLCELL_X32 FILLER_8_317 ();
 FILLCELL_X16 FILLER_8_349 ();
 FILLCELL_X2 FILLER_8_365 ();
 FILLCELL_X32 FILLER_8_368 ();
 FILLCELL_X16 FILLER_8_400 ();
 FILLCELL_X4 FILLER_8_416 ();
 FILLCELL_X1 FILLER_8_420 ();
 FILLCELL_X4 FILLER_9_1 ();
 FILLCELL_X4 FILLER_9_8 ();
 FILLCELL_X32 FILLER_9_15 ();
 FILLCELL_X32 FILLER_9_47 ();
 FILLCELL_X32 FILLER_9_79 ();
 FILLCELL_X32 FILLER_9_111 ();
 FILLCELL_X4 FILLER_9_143 ();
 FILLCELL_X32 FILLER_9_148 ();
 FILLCELL_X32 FILLER_9_180 ();
 FILLCELL_X32 FILLER_9_212 ();
 FILLCELL_X32 FILLER_9_244 ();
 FILLCELL_X16 FILLER_9_276 ();
 FILLCELL_X2 FILLER_9_292 ();
 FILLCELL_X32 FILLER_9_295 ();
 FILLCELL_X32 FILLER_9_327 ();
 FILLCELL_X32 FILLER_9_359 ();
 FILLCELL_X16 FILLER_9_391 ();
 FILLCELL_X8 FILLER_9_407 ();
 FILLCELL_X4 FILLER_9_415 ();
 FILLCELL_X2 FILLER_9_419 ();
 FILLCELL_X4 FILLER_10_1 ();
 FILLCELL_X2 FILLER_10_8 ();
 FILLCELL_X4 FILLER_10_13 ();
 FILLCELL_X32 FILLER_10_20 ();
 FILLCELL_X16 FILLER_10_52 ();
 FILLCELL_X4 FILLER_10_68 ();
 FILLCELL_X1 FILLER_10_72 ();
 FILLCELL_X32 FILLER_10_74 ();
 FILLCELL_X32 FILLER_10_106 ();
 FILLCELL_X32 FILLER_10_138 ();
 FILLCELL_X32 FILLER_10_170 ();
 FILLCELL_X16 FILLER_10_202 ();
 FILLCELL_X2 FILLER_10_218 ();
 FILLCELL_X32 FILLER_10_221 ();
 FILLCELL_X32 FILLER_10_253 ();
 FILLCELL_X32 FILLER_10_285 ();
 FILLCELL_X32 FILLER_10_317 ();
 FILLCELL_X16 FILLER_10_349 ();
 FILLCELL_X2 FILLER_10_365 ();
 FILLCELL_X32 FILLER_10_368 ();
 FILLCELL_X16 FILLER_10_400 ();
 FILLCELL_X4 FILLER_10_416 ();
 FILLCELL_X1 FILLER_10_420 ();
 FILLCELL_X4 FILLER_11_1 ();
 FILLCELL_X2 FILLER_11_5 ();
 FILLCELL_X2 FILLER_11_10 ();
 FILLCELL_X1 FILLER_11_12 ();
 FILLCELL_X2 FILLER_11_18 ();
 FILLCELL_X32 FILLER_11_29 ();
 FILLCELL_X32 FILLER_11_61 ();
 FILLCELL_X32 FILLER_11_93 ();
 FILLCELL_X16 FILLER_11_125 ();
 FILLCELL_X4 FILLER_11_141 ();
 FILLCELL_X2 FILLER_11_145 ();
 FILLCELL_X32 FILLER_11_148 ();
 FILLCELL_X32 FILLER_11_180 ();
 FILLCELL_X32 FILLER_11_212 ();
 FILLCELL_X32 FILLER_11_244 ();
 FILLCELL_X16 FILLER_11_276 ();
 FILLCELL_X2 FILLER_11_292 ();
 FILLCELL_X32 FILLER_11_295 ();
 FILLCELL_X32 FILLER_11_327 ();
 FILLCELL_X32 FILLER_11_359 ();
 FILLCELL_X16 FILLER_11_391 ();
 FILLCELL_X8 FILLER_11_407 ();
 FILLCELL_X4 FILLER_11_415 ();
 FILLCELL_X2 FILLER_11_419 ();
 FILLCELL_X4 FILLER_12_1 ();
 FILLCELL_X2 FILLER_12_5 ();
 FILLCELL_X2 FILLER_12_10 ();
 FILLCELL_X4 FILLER_12_15 ();
 FILLCELL_X1 FILLER_12_19 ();
 FILLCELL_X2 FILLER_12_23 ();
 FILLCELL_X2 FILLER_12_28 ();
 FILLCELL_X2 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_38 ();
 FILLCELL_X2 FILLER_12_70 ();
 FILLCELL_X1 FILLER_12_72 ();
 FILLCELL_X32 FILLER_12_74 ();
 FILLCELL_X32 FILLER_12_106 ();
 FILLCELL_X32 FILLER_12_138 ();
 FILLCELL_X32 FILLER_12_170 ();
 FILLCELL_X16 FILLER_12_202 ();
 FILLCELL_X2 FILLER_12_218 ();
 FILLCELL_X32 FILLER_12_221 ();
 FILLCELL_X32 FILLER_12_253 ();
 FILLCELL_X32 FILLER_12_285 ();
 FILLCELL_X32 FILLER_12_317 ();
 FILLCELL_X16 FILLER_12_349 ();
 FILLCELL_X2 FILLER_12_365 ();
 FILLCELL_X32 FILLER_12_368 ();
 FILLCELL_X16 FILLER_12_400 ();
 FILLCELL_X4 FILLER_12_416 ();
 FILLCELL_X1 FILLER_12_420 ();
 FILLCELL_X2 FILLER_13_1 ();
 FILLCELL_X2 FILLER_13_6 ();
 FILLCELL_X2 FILLER_13_11 ();
 FILLCELL_X4 FILLER_13_16 ();
 FILLCELL_X2 FILLER_13_20 ();
 FILLCELL_X2 FILLER_13_27 ();
 FILLCELL_X2 FILLER_13_32 ();
 FILLCELL_X1 FILLER_13_34 ();
 FILLCELL_X2 FILLER_13_38 ();
 FILLCELL_X32 FILLER_13_49 ();
 FILLCELL_X32 FILLER_13_81 ();
 FILLCELL_X32 FILLER_13_113 ();
 FILLCELL_X2 FILLER_13_145 ();
 FILLCELL_X32 FILLER_13_148 ();
 FILLCELL_X32 FILLER_13_180 ();
 FILLCELL_X32 FILLER_13_212 ();
 FILLCELL_X32 FILLER_13_244 ();
 FILLCELL_X16 FILLER_13_276 ();
 FILLCELL_X2 FILLER_13_292 ();
 FILLCELL_X32 FILLER_13_295 ();
 FILLCELL_X32 FILLER_13_327 ();
 FILLCELL_X32 FILLER_13_359 ();
 FILLCELL_X16 FILLER_13_391 ();
 FILLCELL_X8 FILLER_13_407 ();
 FILLCELL_X4 FILLER_13_415 ();
 FILLCELL_X2 FILLER_13_419 ();
 FILLCELL_X2 FILLER_14_1 ();
 FILLCELL_X1 FILLER_14_3 ();
 FILLCELL_X2 FILLER_14_7 ();
 FILLCELL_X4 FILLER_14_12 ();
 FILLCELL_X2 FILLER_14_16 ();
 FILLCELL_X4 FILLER_14_21 ();
 FILLCELL_X2 FILLER_14_28 ();
 FILLCELL_X2 FILLER_14_32 ();
 FILLCELL_X2 FILLER_14_43 ();
 FILLCELL_X2 FILLER_14_48 ();
 FILLCELL_X2 FILLER_14_53 ();
 FILLCELL_X4 FILLER_14_58 ();
 FILLCELL_X2 FILLER_14_62 ();
 FILLCELL_X4 FILLER_14_67 ();
 FILLCELL_X2 FILLER_14_71 ();
 FILLCELL_X32 FILLER_14_74 ();
 FILLCELL_X32 FILLER_14_106 ();
 FILLCELL_X32 FILLER_14_138 ();
 FILLCELL_X32 FILLER_14_170 ();
 FILLCELL_X16 FILLER_14_202 ();
 FILLCELL_X2 FILLER_14_218 ();
 FILLCELL_X32 FILLER_14_221 ();
 FILLCELL_X32 FILLER_14_253 ();
 FILLCELL_X32 FILLER_14_285 ();
 FILLCELL_X32 FILLER_14_317 ();
 FILLCELL_X16 FILLER_14_349 ();
 FILLCELL_X2 FILLER_14_365 ();
 FILLCELL_X32 FILLER_14_368 ();
 FILLCELL_X16 FILLER_14_400 ();
 FILLCELL_X4 FILLER_14_416 ();
 FILLCELL_X1 FILLER_14_420 ();
 FILLCELL_X2 FILLER_15_1 ();
 FILLCELL_X1 FILLER_15_3 ();
 FILLCELL_X2 FILLER_15_21 ();
 FILLCELL_X4 FILLER_15_26 ();
 FILLCELL_X2 FILLER_15_34 ();
 FILLCELL_X2 FILLER_15_53 ();
 FILLCELL_X4 FILLER_15_60 ();
 FILLCELL_X1 FILLER_15_64 ();
 FILLCELL_X2 FILLER_15_82 ();
 FILLCELL_X4 FILLER_15_87 ();
 FILLCELL_X2 FILLER_15_91 ();
 FILLCELL_X32 FILLER_15_96 ();
 FILLCELL_X16 FILLER_15_128 ();
 FILLCELL_X2 FILLER_15_144 ();
 FILLCELL_X1 FILLER_15_146 ();
 FILLCELL_X32 FILLER_15_148 ();
 FILLCELL_X32 FILLER_15_180 ();
 FILLCELL_X32 FILLER_15_212 ();
 FILLCELL_X32 FILLER_15_244 ();
 FILLCELL_X16 FILLER_15_276 ();
 FILLCELL_X2 FILLER_15_292 ();
 FILLCELL_X32 FILLER_15_295 ();
 FILLCELL_X32 FILLER_15_327 ();
 FILLCELL_X32 FILLER_15_359 ();
 FILLCELL_X16 FILLER_15_391 ();
 FILLCELL_X8 FILLER_15_407 ();
 FILLCELL_X4 FILLER_15_415 ();
 FILLCELL_X2 FILLER_15_419 ();
 FILLCELL_X2 FILLER_16_1 ();
 FILLCELL_X2 FILLER_16_20 ();
 FILLCELL_X1 FILLER_16_22 ();
 FILLCELL_X2 FILLER_16_29 ();
 FILLCELL_X2 FILLER_16_40 ();
 FILLCELL_X2 FILLER_16_51 ();
 FILLCELL_X2 FILLER_16_70 ();
 FILLCELL_X1 FILLER_16_72 ();
 FILLCELL_X2 FILLER_16_74 ();
 FILLCELL_X1 FILLER_16_76 ();
 FILLCELL_X2 FILLER_16_94 ();
 FILLCELL_X2 FILLER_16_99 ();
 FILLCELL_X32 FILLER_16_106 ();
 FILLCELL_X32 FILLER_16_138 ();
 FILLCELL_X32 FILLER_16_170 ();
 FILLCELL_X16 FILLER_16_202 ();
 FILLCELL_X2 FILLER_16_218 ();
 FILLCELL_X32 FILLER_16_221 ();
 FILLCELL_X32 FILLER_16_253 ();
 FILLCELL_X32 FILLER_16_285 ();
 FILLCELL_X32 FILLER_16_317 ();
 FILLCELL_X16 FILLER_16_349 ();
 FILLCELL_X2 FILLER_16_365 ();
 FILLCELL_X32 FILLER_16_368 ();
 FILLCELL_X16 FILLER_16_400 ();
 FILLCELL_X4 FILLER_16_416 ();
 FILLCELL_X1 FILLER_16_420 ();
 FILLCELL_X4 FILLER_17_1 ();
 FILLCELL_X1 FILLER_17_5 ();
 FILLCELL_X2 FILLER_17_9 ();
 FILLCELL_X1 FILLER_17_11 ();
 FILLCELL_X2 FILLER_17_15 ();
 FILLCELL_X2 FILLER_17_20 ();
 FILLCELL_X2 FILLER_17_25 ();
 FILLCELL_X1 FILLER_17_27 ();
 FILLCELL_X2 FILLER_17_37 ();
 FILLCELL_X2 FILLER_17_48 ();
 FILLCELL_X4 FILLER_17_53 ();
 FILLCELL_X2 FILLER_17_61 ();
 FILLCELL_X2 FILLER_17_65 ();
 FILLCELL_X4 FILLER_17_71 ();
 FILLCELL_X1 FILLER_17_75 ();
 FILLCELL_X2 FILLER_17_79 ();
 FILLCELL_X2 FILLER_17_94 ();
 FILLCELL_X2 FILLER_17_106 ();
 FILLCELL_X32 FILLER_17_113 ();
 FILLCELL_X2 FILLER_17_145 ();
 FILLCELL_X32 FILLER_17_148 ();
 FILLCELL_X32 FILLER_17_180 ();
 FILLCELL_X32 FILLER_17_212 ();
 FILLCELL_X32 FILLER_17_244 ();
 FILLCELL_X16 FILLER_17_276 ();
 FILLCELL_X2 FILLER_17_292 ();
 FILLCELL_X32 FILLER_17_295 ();
 FILLCELL_X32 FILLER_17_327 ();
 FILLCELL_X32 FILLER_17_359 ();
 FILLCELL_X16 FILLER_17_391 ();
 FILLCELL_X8 FILLER_17_407 ();
 FILLCELL_X4 FILLER_17_415 ();
 FILLCELL_X2 FILLER_17_419 ();
 FILLCELL_X4 FILLER_18_1 ();
 FILLCELL_X2 FILLER_18_5 ();
 FILLCELL_X2 FILLER_18_10 ();
 FILLCELL_X2 FILLER_18_19 ();
 FILLCELL_X2 FILLER_18_25 ();
 FILLCELL_X1 FILLER_18_27 ();
 FILLCELL_X2 FILLER_18_31 ();
 FILLCELL_X2 FILLER_18_39 ();
 FILLCELL_X2 FILLER_18_45 ();
 FILLCELL_X1 FILLER_18_47 ();
 FILLCELL_X2 FILLER_18_51 ();
 FILLCELL_X2 FILLER_18_59 ();
 FILLCELL_X2 FILLER_18_71 ();
 FILLCELL_X2 FILLER_18_74 ();
 FILLCELL_X2 FILLER_18_78 ();
 FILLCELL_X2 FILLER_18_84 ();
 FILLCELL_X1 FILLER_18_86 ();
 FILLCELL_X4 FILLER_18_100 ();
 FILLCELL_X1 FILLER_18_104 ();
 FILLCELL_X32 FILLER_18_114 ();
 FILLCELL_X32 FILLER_18_146 ();
 FILLCELL_X32 FILLER_18_178 ();
 FILLCELL_X8 FILLER_18_210 ();
 FILLCELL_X2 FILLER_18_218 ();
 FILLCELL_X32 FILLER_18_221 ();
 FILLCELL_X32 FILLER_18_253 ();
 FILLCELL_X32 FILLER_18_285 ();
 FILLCELL_X32 FILLER_18_317 ();
 FILLCELL_X16 FILLER_18_349 ();
 FILLCELL_X2 FILLER_18_365 ();
 FILLCELL_X32 FILLER_18_368 ();
 FILLCELL_X16 FILLER_18_400 ();
 FILLCELL_X4 FILLER_18_416 ();
 FILLCELL_X1 FILLER_18_420 ();
 FILLCELL_X2 FILLER_19_1 ();
 FILLCELL_X2 FILLER_19_20 ();
 FILLCELL_X2 FILLER_19_24 ();
 FILLCELL_X2 FILLER_19_30 ();
 FILLCELL_X1 FILLER_19_32 ();
 FILLCELL_X2 FILLER_19_38 ();
 FILLCELL_X2 FILLER_19_44 ();
 FILLCELL_X2 FILLER_19_51 ();
 FILLCELL_X4 FILLER_19_58 ();
 FILLCELL_X4 FILLER_19_65 ();
 FILLCELL_X2 FILLER_19_73 ();
 FILLCELL_X2 FILLER_19_77 ();
 FILLCELL_X2 FILLER_19_83 ();
 FILLCELL_X2 FILLER_19_94 ();
 FILLCELL_X2 FILLER_19_109 ();
 FILLCELL_X2 FILLER_19_120 ();
 FILLCELL_X16 FILLER_19_131 ();
 FILLCELL_X32 FILLER_19_148 ();
 FILLCELL_X32 FILLER_19_180 ();
 FILLCELL_X32 FILLER_19_212 ();
 FILLCELL_X32 FILLER_19_244 ();
 FILLCELL_X16 FILLER_19_276 ();
 FILLCELL_X2 FILLER_19_292 ();
 FILLCELL_X32 FILLER_19_295 ();
 FILLCELL_X32 FILLER_19_327 ();
 FILLCELL_X32 FILLER_19_359 ();
 FILLCELL_X16 FILLER_19_391 ();
 FILLCELL_X8 FILLER_19_407 ();
 FILLCELL_X4 FILLER_19_415 ();
 FILLCELL_X2 FILLER_19_419 ();
 FILLCELL_X2 FILLER_20_1 ();
 FILLCELL_X1 FILLER_20_3 ();
 FILLCELL_X2 FILLER_20_7 ();
 FILLCELL_X2 FILLER_20_13 ();
 FILLCELL_X2 FILLER_20_19 ();
 FILLCELL_X1 FILLER_20_21 ();
 FILLCELL_X2 FILLER_20_25 ();
 FILLCELL_X4 FILLER_20_31 ();
 FILLCELL_X1 FILLER_20_35 ();
 FILLCELL_X2 FILLER_20_39 ();
 FILLCELL_X2 FILLER_20_44 ();
 FILLCELL_X2 FILLER_20_49 ();
 FILLCELL_X2 FILLER_20_55 ();
 FILLCELL_X1 FILLER_20_57 ();
 FILLCELL_X2 FILLER_20_61 ();
 FILLCELL_X2 FILLER_20_66 ();
 FILLCELL_X2 FILLER_20_71 ();
 FILLCELL_X2 FILLER_20_74 ();
 FILLCELL_X2 FILLER_20_85 ();
 FILLCELL_X4 FILLER_20_93 ();
 FILLCELL_X1 FILLER_20_97 ();
 FILLCELL_X2 FILLER_20_107 ();
 FILLCELL_X2 FILLER_20_118 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X16 FILLER_20_193 ();
 FILLCELL_X8 FILLER_20_209 ();
 FILLCELL_X2 FILLER_20_217 ();
 FILLCELL_X1 FILLER_20_219 ();
 FILLCELL_X32 FILLER_20_221 ();
 FILLCELL_X32 FILLER_20_253 ();
 FILLCELL_X32 FILLER_20_285 ();
 FILLCELL_X32 FILLER_20_317 ();
 FILLCELL_X16 FILLER_20_349 ();
 FILLCELL_X2 FILLER_20_365 ();
 FILLCELL_X32 FILLER_20_368 ();
 FILLCELL_X16 FILLER_20_400 ();
 FILLCELL_X4 FILLER_20_416 ();
 FILLCELL_X1 FILLER_20_420 ();
 FILLCELL_X4 FILLER_21_1 ();
 FILLCELL_X1 FILLER_21_5 ();
 FILLCELL_X2 FILLER_21_9 ();
 FILLCELL_X2 FILLER_21_14 ();
 FILLCELL_X1 FILLER_21_16 ();
 FILLCELL_X2 FILLER_21_20 ();
 FILLCELL_X4 FILLER_21_27 ();
 FILLCELL_X2 FILLER_21_31 ();
 FILLCELL_X2 FILLER_21_46 ();
 FILLCELL_X1 FILLER_21_48 ();
 FILLCELL_X4 FILLER_21_66 ();
 FILLCELL_X1 FILLER_21_70 ();
 FILLCELL_X2 FILLER_21_74 ();
 FILLCELL_X2 FILLER_21_79 ();
 FILLCELL_X2 FILLER_21_85 ();
 FILLCELL_X2 FILLER_21_94 ();
 FILLCELL_X2 FILLER_21_106 ();
 FILLCELL_X2 FILLER_21_111 ();
 FILLCELL_X2 FILLER_21_116 ();
 FILLCELL_X16 FILLER_21_121 ();
 FILLCELL_X8 FILLER_21_137 ();
 FILLCELL_X2 FILLER_21_145 ();
 FILLCELL_X32 FILLER_21_148 ();
 FILLCELL_X32 FILLER_21_180 ();
 FILLCELL_X32 FILLER_21_212 ();
 FILLCELL_X32 FILLER_21_244 ();
 FILLCELL_X16 FILLER_21_276 ();
 FILLCELL_X2 FILLER_21_292 ();
 FILLCELL_X32 FILLER_21_295 ();
 FILLCELL_X32 FILLER_21_327 ();
 FILLCELL_X32 FILLER_21_359 ();
 FILLCELL_X16 FILLER_21_391 ();
 FILLCELL_X8 FILLER_21_407 ();
 FILLCELL_X4 FILLER_21_415 ();
 FILLCELL_X2 FILLER_21_419 ();
 FILLCELL_X4 FILLER_22_1 ();
 FILLCELL_X2 FILLER_22_5 ();
 FILLCELL_X2 FILLER_22_14 ();
 FILLCELL_X2 FILLER_22_23 ();
 FILLCELL_X2 FILLER_22_27 ();
 FILLCELL_X2 FILLER_22_46 ();
 FILLCELL_X2 FILLER_22_51 ();
 FILLCELL_X2 FILLER_22_60 ();
 FILLCELL_X4 FILLER_22_67 ();
 FILLCELL_X2 FILLER_22_71 ();
 FILLCELL_X2 FILLER_22_74 ();
 FILLCELL_X1 FILLER_22_76 ();
 FILLCELL_X2 FILLER_22_84 ();
 FILLCELL_X4 FILLER_22_93 ();
 FILLCELL_X2 FILLER_22_107 ();
 FILLCELL_X32 FILLER_22_126 ();
 FILLCELL_X32 FILLER_22_158 ();
 FILLCELL_X16 FILLER_22_190 ();
 FILLCELL_X8 FILLER_22_206 ();
 FILLCELL_X4 FILLER_22_214 ();
 FILLCELL_X2 FILLER_22_218 ();
 FILLCELL_X32 FILLER_22_221 ();
 FILLCELL_X32 FILLER_22_253 ();
 FILLCELL_X32 FILLER_22_285 ();
 FILLCELL_X32 FILLER_22_317 ();
 FILLCELL_X16 FILLER_22_349 ();
 FILLCELL_X2 FILLER_22_365 ();
 FILLCELL_X32 FILLER_22_368 ();
 FILLCELL_X16 FILLER_22_400 ();
 FILLCELL_X4 FILLER_22_416 ();
 FILLCELL_X1 FILLER_22_420 ();
 FILLCELL_X2 FILLER_23_1 ();
 FILLCELL_X4 FILLER_23_20 ();
 FILLCELL_X1 FILLER_23_24 ();
 FILLCELL_X2 FILLER_23_31 ();
 FILLCELL_X2 FILLER_23_39 ();
 FILLCELL_X2 FILLER_23_48 ();
 FILLCELL_X4 FILLER_23_55 ();
 FILLCELL_X2 FILLER_23_59 ();
 FILLCELL_X2 FILLER_23_65 ();
 FILLCELL_X8 FILLER_23_84 ();
 FILLCELL_X1 FILLER_23_92 ();
 FILLCELL_X2 FILLER_23_100 ();
 FILLCELL_X2 FILLER_23_112 ();
 FILLCELL_X1 FILLER_23_114 ();
 FILLCELL_X8 FILLER_23_132 ();
 FILLCELL_X4 FILLER_23_140 ();
 FILLCELL_X2 FILLER_23_144 ();
 FILLCELL_X1 FILLER_23_146 ();
 FILLCELL_X32 FILLER_23_148 ();
 FILLCELL_X32 FILLER_23_180 ();
 FILLCELL_X32 FILLER_23_212 ();
 FILLCELL_X32 FILLER_23_244 ();
 FILLCELL_X16 FILLER_23_276 ();
 FILLCELL_X2 FILLER_23_292 ();
 FILLCELL_X32 FILLER_23_295 ();
 FILLCELL_X32 FILLER_23_327 ();
 FILLCELL_X32 FILLER_23_359 ();
 FILLCELL_X16 FILLER_23_391 ();
 FILLCELL_X8 FILLER_23_407 ();
 FILLCELL_X4 FILLER_23_415 ();
 FILLCELL_X2 FILLER_23_419 ();
 FILLCELL_X4 FILLER_24_1 ();
 FILLCELL_X1 FILLER_24_5 ();
 FILLCELL_X2 FILLER_24_9 ();
 FILLCELL_X4 FILLER_24_15 ();
 FILLCELL_X2 FILLER_24_22 ();
 FILLCELL_X4 FILLER_24_29 ();
 FILLCELL_X1 FILLER_24_33 ();
 FILLCELL_X2 FILLER_24_37 ();
 FILLCELL_X4 FILLER_24_42 ();
 FILLCELL_X2 FILLER_24_46 ();
 FILLCELL_X2 FILLER_24_65 ();
 FILLCELL_X2 FILLER_24_71 ();
 FILLCELL_X4 FILLER_24_74 ();
 FILLCELL_X2 FILLER_24_78 ();
 FILLCELL_X2 FILLER_24_85 ();
 FILLCELL_X4 FILLER_24_91 ();
 FILLCELL_X1 FILLER_24_95 ();
 FILLCELL_X2 FILLER_24_100 ();
 FILLCELL_X1 FILLER_24_102 ();
 FILLCELL_X2 FILLER_24_106 ();
 FILLCELL_X2 FILLER_24_113 ();
 FILLCELL_X32 FILLER_24_118 ();
 FILLCELL_X32 FILLER_24_150 ();
 FILLCELL_X32 FILLER_24_182 ();
 FILLCELL_X4 FILLER_24_214 ();
 FILLCELL_X2 FILLER_24_218 ();
 FILLCELL_X32 FILLER_24_221 ();
 FILLCELL_X32 FILLER_24_253 ();
 FILLCELL_X32 FILLER_24_285 ();
 FILLCELL_X32 FILLER_24_317 ();
 FILLCELL_X16 FILLER_24_349 ();
 FILLCELL_X2 FILLER_24_365 ();
 FILLCELL_X32 FILLER_24_368 ();
 FILLCELL_X16 FILLER_24_400 ();
 FILLCELL_X4 FILLER_24_416 ();
 FILLCELL_X1 FILLER_24_420 ();
 FILLCELL_X2 FILLER_25_1 ();
 FILLCELL_X4 FILLER_25_6 ();
 FILLCELL_X1 FILLER_25_10 ();
 FILLCELL_X4 FILLER_25_15 ();
 FILLCELL_X2 FILLER_25_19 ();
 FILLCELL_X2 FILLER_25_27 ();
 FILLCELL_X2 FILLER_25_33 ();
 FILLCELL_X2 FILLER_25_37 ();
 FILLCELL_X2 FILLER_25_42 ();
 FILLCELL_X2 FILLER_25_51 ();
 FILLCELL_X2 FILLER_25_57 ();
 FILLCELL_X2 FILLER_25_61 ();
 FILLCELL_X2 FILLER_25_66 ();
 FILLCELL_X4 FILLER_25_71 ();
 FILLCELL_X2 FILLER_25_75 ();
 FILLCELL_X2 FILLER_25_80 ();
 FILLCELL_X4 FILLER_25_85 ();
 FILLCELL_X2 FILLER_25_92 ();
 FILLCELL_X2 FILLER_25_98 ();
 FILLCELL_X2 FILLER_25_103 ();
 FILLCELL_X2 FILLER_25_115 ();
 FILLCELL_X8 FILLER_25_134 ();
 FILLCELL_X4 FILLER_25_142 ();
 FILLCELL_X1 FILLER_25_146 ();
 FILLCELL_X32 FILLER_25_148 ();
 FILLCELL_X32 FILLER_25_180 ();
 FILLCELL_X32 FILLER_25_212 ();
 FILLCELL_X32 FILLER_25_244 ();
 FILLCELL_X16 FILLER_25_276 ();
 FILLCELL_X2 FILLER_25_292 ();
 FILLCELL_X32 FILLER_25_295 ();
 FILLCELL_X32 FILLER_25_327 ();
 FILLCELL_X32 FILLER_25_359 ();
 FILLCELL_X16 FILLER_25_391 ();
 FILLCELL_X8 FILLER_25_407 ();
 FILLCELL_X4 FILLER_25_415 ();
 FILLCELL_X2 FILLER_25_419 ();
 FILLCELL_X2 FILLER_26_1 ();
 FILLCELL_X4 FILLER_26_20 ();
 FILLCELL_X1 FILLER_26_24 ();
 FILLCELL_X2 FILLER_26_42 ();
 FILLCELL_X4 FILLER_26_51 ();
 FILLCELL_X2 FILLER_26_59 ();
 FILLCELL_X2 FILLER_26_64 ();
 FILLCELL_X1 FILLER_26_66 ();
 FILLCELL_X2 FILLER_26_71 ();
 FILLCELL_X4 FILLER_26_74 ();
 FILLCELL_X2 FILLER_26_78 ();
 FILLCELL_X2 FILLER_26_83 ();
 FILLCELL_X1 FILLER_26_85 ();
 FILLCELL_X4 FILLER_26_91 ();
 FILLCELL_X2 FILLER_26_95 ();
 FILLCELL_X4 FILLER_26_114 ();
 FILLCELL_X1 FILLER_26_118 ();
 FILLCELL_X2 FILLER_26_124 ();
 FILLCELL_X2 FILLER_26_136 ();
 FILLCELL_X32 FILLER_26_141 ();
 FILLCELL_X32 FILLER_26_173 ();
 FILLCELL_X8 FILLER_26_205 ();
 FILLCELL_X4 FILLER_26_213 ();
 FILLCELL_X2 FILLER_26_217 ();
 FILLCELL_X1 FILLER_26_219 ();
 FILLCELL_X32 FILLER_26_221 ();
 FILLCELL_X32 FILLER_26_253 ();
 FILLCELL_X32 FILLER_26_285 ();
 FILLCELL_X32 FILLER_26_317 ();
 FILLCELL_X16 FILLER_26_349 ();
 FILLCELL_X2 FILLER_26_365 ();
 FILLCELL_X32 FILLER_26_368 ();
 FILLCELL_X16 FILLER_26_400 ();
 FILLCELL_X4 FILLER_26_416 ();
 FILLCELL_X1 FILLER_26_420 ();
 FILLCELL_X4 FILLER_27_1 ();
 FILLCELL_X2 FILLER_27_5 ();
 FILLCELL_X2 FILLER_27_10 ();
 FILLCELL_X2 FILLER_27_19 ();
 FILLCELL_X2 FILLER_27_24 ();
 FILLCELL_X4 FILLER_27_30 ();
 FILLCELL_X1 FILLER_27_34 ();
 FILLCELL_X2 FILLER_27_38 ();
 FILLCELL_X2 FILLER_27_43 ();
 FILLCELL_X2 FILLER_27_50 ();
 FILLCELL_X2 FILLER_27_69 ();
 FILLCELL_X2 FILLER_27_73 ();
 FILLCELL_X2 FILLER_27_79 ();
 FILLCELL_X2 FILLER_27_86 ();
 FILLCELL_X4 FILLER_27_92 ();
 FILLCELL_X2 FILLER_27_100 ();
 FILLCELL_X2 FILLER_27_105 ();
 FILLCELL_X1 FILLER_27_107 ();
 FILLCELL_X4 FILLER_27_110 ();
 FILLCELL_X2 FILLER_27_114 ();
 FILLCELL_X2 FILLER_27_122 ();
 FILLCELL_X8 FILLER_27_134 ();
 FILLCELL_X4 FILLER_27_142 ();
 FILLCELL_X1 FILLER_27_146 ();
 FILLCELL_X32 FILLER_27_148 ();
 FILLCELL_X32 FILLER_27_180 ();
 FILLCELL_X32 FILLER_27_212 ();
 FILLCELL_X32 FILLER_27_244 ();
 FILLCELL_X16 FILLER_27_276 ();
 FILLCELL_X2 FILLER_27_292 ();
 FILLCELL_X32 FILLER_27_295 ();
 FILLCELL_X32 FILLER_27_327 ();
 FILLCELL_X32 FILLER_27_359 ();
 FILLCELL_X16 FILLER_27_391 ();
 FILLCELL_X8 FILLER_27_407 ();
 FILLCELL_X4 FILLER_27_415 ();
 FILLCELL_X2 FILLER_27_419 ();
 FILLCELL_X2 FILLER_28_1 ();
 FILLCELL_X1 FILLER_28_3 ();
 FILLCELL_X4 FILLER_28_7 ();
 FILLCELL_X1 FILLER_28_11 ();
 FILLCELL_X4 FILLER_28_16 ();
 FILLCELL_X4 FILLER_28_24 ();
 FILLCELL_X2 FILLER_28_28 ();
 FILLCELL_X2 FILLER_28_34 ();
 FILLCELL_X2 FILLER_28_40 ();
 FILLCELL_X1 FILLER_28_42 ();
 FILLCELL_X2 FILLER_28_46 ();
 FILLCELL_X4 FILLER_28_53 ();
 FILLCELL_X2 FILLER_28_57 ();
 FILLCELL_X2 FILLER_28_62 ();
 FILLCELL_X2 FILLER_28_71 ();
 FILLCELL_X4 FILLER_28_74 ();
 FILLCELL_X1 FILLER_28_78 ();
 FILLCELL_X2 FILLER_28_86 ();
 FILLCELL_X2 FILLER_28_92 ();
 FILLCELL_X2 FILLER_28_97 ();
 FILLCELL_X2 FILLER_28_116 ();
 FILLCELL_X2 FILLER_28_121 ();
 FILLCELL_X2 FILLER_28_136 ();
 FILLCELL_X32 FILLER_28_142 ();
 FILLCELL_X32 FILLER_28_174 ();
 FILLCELL_X8 FILLER_28_206 ();
 FILLCELL_X4 FILLER_28_214 ();
 FILLCELL_X2 FILLER_28_218 ();
 FILLCELL_X32 FILLER_28_221 ();
 FILLCELL_X32 FILLER_28_253 ();
 FILLCELL_X32 FILLER_28_285 ();
 FILLCELL_X32 FILLER_28_317 ();
 FILLCELL_X16 FILLER_28_349 ();
 FILLCELL_X2 FILLER_28_365 ();
 FILLCELL_X32 FILLER_28_368 ();
 FILLCELL_X16 FILLER_28_400 ();
 FILLCELL_X4 FILLER_28_416 ();
 FILLCELL_X1 FILLER_28_420 ();
 FILLCELL_X4 FILLER_29_1 ();
 FILLCELL_X1 FILLER_29_5 ();
 FILLCELL_X4 FILLER_29_23 ();
 FILLCELL_X2 FILLER_29_44 ();
 FILLCELL_X2 FILLER_29_49 ();
 FILLCELL_X2 FILLER_29_61 ();
 FILLCELL_X2 FILLER_29_67 ();
 FILLCELL_X2 FILLER_29_72 ();
 FILLCELL_X2 FILLER_29_76 ();
 FILLCELL_X2 FILLER_29_81 ();
 FILLCELL_X4 FILLER_29_87 ();
 FILLCELL_X2 FILLER_29_91 ();
 FILLCELL_X4 FILLER_29_110 ();
 FILLCELL_X2 FILLER_29_117 ();
 FILLCELL_X2 FILLER_29_129 ();
 FILLCELL_X8 FILLER_29_134 ();
 FILLCELL_X4 FILLER_29_142 ();
 FILLCELL_X1 FILLER_29_146 ();
 FILLCELL_X32 FILLER_29_148 ();
 FILLCELL_X32 FILLER_29_180 ();
 FILLCELL_X32 FILLER_29_212 ();
 FILLCELL_X32 FILLER_29_244 ();
 FILLCELL_X16 FILLER_29_276 ();
 FILLCELL_X2 FILLER_29_292 ();
 FILLCELL_X32 FILLER_29_295 ();
 FILLCELL_X32 FILLER_29_327 ();
 FILLCELL_X32 FILLER_29_359 ();
 FILLCELL_X16 FILLER_29_391 ();
 FILLCELL_X8 FILLER_29_407 ();
 FILLCELL_X4 FILLER_29_415 ();
 FILLCELL_X2 FILLER_29_419 ();
 FILLCELL_X2 FILLER_30_1 ();
 FILLCELL_X1 FILLER_30_3 ();
 FILLCELL_X2 FILLER_30_7 ();
 FILLCELL_X2 FILLER_30_12 ();
 FILLCELL_X2 FILLER_30_17 ();
 FILLCELL_X2 FILLER_30_22 ();
 FILLCELL_X2 FILLER_30_33 ();
 FILLCELL_X2 FILLER_30_38 ();
 FILLCELL_X2 FILLER_30_46 ();
 FILLCELL_X2 FILLER_30_55 ();
 FILLCELL_X2 FILLER_30_66 ();
 FILLCELL_X2 FILLER_30_71 ();
 FILLCELL_X4 FILLER_30_74 ();
 FILLCELL_X4 FILLER_30_81 ();
 FILLCELL_X1 FILLER_30_85 ();
 FILLCELL_X2 FILLER_30_90 ();
 FILLCELL_X1 FILLER_30_92 ();
 FILLCELL_X2 FILLER_30_96 ();
 FILLCELL_X2 FILLER_30_101 ();
 FILLCELL_X1 FILLER_30_103 ();
 FILLCELL_X2 FILLER_30_121 ();
 FILLCELL_X32 FILLER_30_126 ();
 FILLCELL_X32 FILLER_30_158 ();
 FILLCELL_X16 FILLER_30_190 ();
 FILLCELL_X8 FILLER_30_206 ();
 FILLCELL_X4 FILLER_30_214 ();
 FILLCELL_X2 FILLER_30_218 ();
 FILLCELL_X32 FILLER_30_221 ();
 FILLCELL_X32 FILLER_30_253 ();
 FILLCELL_X32 FILLER_30_285 ();
 FILLCELL_X32 FILLER_30_317 ();
 FILLCELL_X16 FILLER_30_349 ();
 FILLCELL_X2 FILLER_30_365 ();
 FILLCELL_X32 FILLER_30_368 ();
 FILLCELL_X16 FILLER_30_400 ();
 FILLCELL_X4 FILLER_30_416 ();
 FILLCELL_X1 FILLER_30_420 ();
 FILLCELL_X4 FILLER_31_1 ();
 FILLCELL_X2 FILLER_31_8 ();
 FILLCELL_X2 FILLER_31_13 ();
 FILLCELL_X4 FILLER_31_19 ();
 FILLCELL_X2 FILLER_31_27 ();
 FILLCELL_X2 FILLER_31_32 ();
 FILLCELL_X2 FILLER_31_38 ();
 FILLCELL_X1 FILLER_31_40 ();
 FILLCELL_X2 FILLER_31_46 ();
 FILLCELL_X2 FILLER_31_53 ();
 FILLCELL_X4 FILLER_31_64 ();
 FILLCELL_X2 FILLER_31_71 ();
 FILLCELL_X2 FILLER_31_77 ();
 FILLCELL_X2 FILLER_31_92 ();
 FILLCELL_X4 FILLER_31_101 ();
 FILLCELL_X2 FILLER_31_105 ();
 FILLCELL_X2 FILLER_31_117 ();
 FILLCELL_X2 FILLER_31_128 ();
 FILLCELL_X8 FILLER_31_133 ();
 FILLCELL_X4 FILLER_31_141 ();
 FILLCELL_X2 FILLER_31_145 ();
 FILLCELL_X32 FILLER_31_148 ();
 FILLCELL_X32 FILLER_31_180 ();
 FILLCELL_X32 FILLER_31_212 ();
 FILLCELL_X32 FILLER_31_244 ();
 FILLCELL_X16 FILLER_31_276 ();
 FILLCELL_X2 FILLER_31_292 ();
 FILLCELL_X32 FILLER_31_295 ();
 FILLCELL_X32 FILLER_31_327 ();
 FILLCELL_X32 FILLER_31_359 ();
 FILLCELL_X16 FILLER_31_391 ();
 FILLCELL_X8 FILLER_31_407 ();
 FILLCELL_X4 FILLER_31_415 ();
 FILLCELL_X2 FILLER_31_419 ();
 FILLCELL_X2 FILLER_32_1 ();
 FILLCELL_X2 FILLER_32_5 ();
 FILLCELL_X2 FILLER_32_10 ();
 FILLCELL_X2 FILLER_32_29 ();
 FILLCELL_X1 FILLER_32_31 ();
 FILLCELL_X2 FILLER_32_39 ();
 FILLCELL_X2 FILLER_32_50 ();
 FILLCELL_X2 FILLER_32_62 ();
 FILLCELL_X2 FILLER_32_67 ();
 FILLCELL_X2 FILLER_32_71 ();
 FILLCELL_X4 FILLER_32_74 ();
 FILLCELL_X2 FILLER_32_85 ();
 FILLCELL_X1 FILLER_32_87 ();
 FILLCELL_X2 FILLER_32_105 ();
 FILLCELL_X2 FILLER_32_109 ();
 FILLCELL_X2 FILLER_32_114 ();
 FILLCELL_X1 FILLER_32_116 ();
 FILLCELL_X2 FILLER_32_127 ();
 FILLCELL_X32 FILLER_32_138 ();
 FILLCELL_X32 FILLER_32_170 ();
 FILLCELL_X16 FILLER_32_202 ();
 FILLCELL_X2 FILLER_32_218 ();
 FILLCELL_X32 FILLER_32_221 ();
 FILLCELL_X32 FILLER_32_253 ();
 FILLCELL_X32 FILLER_32_285 ();
 FILLCELL_X32 FILLER_32_317 ();
 FILLCELL_X16 FILLER_32_349 ();
 FILLCELL_X2 FILLER_32_365 ();
 FILLCELL_X32 FILLER_32_368 ();
 FILLCELL_X16 FILLER_32_400 ();
 FILLCELL_X4 FILLER_32_416 ();
 FILLCELL_X1 FILLER_32_420 ();
 FILLCELL_X2 FILLER_33_1 ();
 FILLCELL_X2 FILLER_33_5 ();
 FILLCELL_X2 FILLER_33_11 ();
 FILLCELL_X1 FILLER_33_13 ();
 FILLCELL_X2 FILLER_33_17 ();
 FILLCELL_X2 FILLER_33_22 ();
 FILLCELL_X2 FILLER_33_27 ();
 FILLCELL_X2 FILLER_33_33 ();
 FILLCELL_X2 FILLER_33_39 ();
 FILLCELL_X4 FILLER_33_45 ();
 FILLCELL_X2 FILLER_33_52 ();
 FILLCELL_X2 FILLER_33_58 ();
 FILLCELL_X2 FILLER_33_64 ();
 FILLCELL_X1 FILLER_33_66 ();
 FILLCELL_X4 FILLER_33_70 ();
 FILLCELL_X2 FILLER_33_77 ();
 FILLCELL_X2 FILLER_33_84 ();
 FILLCELL_X2 FILLER_33_90 ();
 FILLCELL_X2 FILLER_33_95 ();
 FILLCELL_X2 FILLER_33_106 ();
 FILLCELL_X2 FILLER_33_118 ();
 FILLCELL_X2 FILLER_33_130 ();
 FILLCELL_X8 FILLER_33_135 ();
 FILLCELL_X4 FILLER_33_143 ();
 FILLCELL_X32 FILLER_33_148 ();
 FILLCELL_X32 FILLER_33_180 ();
 FILLCELL_X32 FILLER_33_212 ();
 FILLCELL_X32 FILLER_33_244 ();
 FILLCELL_X16 FILLER_33_276 ();
 FILLCELL_X2 FILLER_33_292 ();
 FILLCELL_X32 FILLER_33_295 ();
 FILLCELL_X32 FILLER_33_327 ();
 FILLCELL_X32 FILLER_33_359 ();
 FILLCELL_X16 FILLER_33_391 ();
 FILLCELL_X8 FILLER_33_407 ();
 FILLCELL_X4 FILLER_33_415 ();
 FILLCELL_X2 FILLER_33_419 ();
 FILLCELL_X2 FILLER_34_1 ();
 FILLCELL_X2 FILLER_34_20 ();
 FILLCELL_X2 FILLER_34_25 ();
 FILLCELL_X2 FILLER_34_30 ();
 FILLCELL_X2 FILLER_34_39 ();
 FILLCELL_X2 FILLER_34_48 ();
 FILLCELL_X4 FILLER_34_55 ();
 FILLCELL_X1 FILLER_34_59 ();
 FILLCELL_X2 FILLER_34_64 ();
 FILLCELL_X2 FILLER_34_70 ();
 FILLCELL_X1 FILLER_34_72 ();
 FILLCELL_X2 FILLER_34_74 ();
 FILLCELL_X2 FILLER_34_83 ();
 FILLCELL_X2 FILLER_34_102 ();
 FILLCELL_X4 FILLER_34_109 ();
 FILLCELL_X1 FILLER_34_113 ();
 FILLCELL_X2 FILLER_34_127 ();
 FILLCELL_X32 FILLER_34_136 ();
 FILLCELL_X32 FILLER_34_168 ();
 FILLCELL_X16 FILLER_34_200 ();
 FILLCELL_X4 FILLER_34_216 ();
 FILLCELL_X32 FILLER_34_221 ();
 FILLCELL_X32 FILLER_34_253 ();
 FILLCELL_X32 FILLER_34_285 ();
 FILLCELL_X32 FILLER_34_317 ();
 FILLCELL_X16 FILLER_34_349 ();
 FILLCELL_X2 FILLER_34_365 ();
 FILLCELL_X32 FILLER_34_368 ();
 FILLCELL_X16 FILLER_34_400 ();
 FILLCELL_X4 FILLER_34_416 ();
 FILLCELL_X1 FILLER_34_420 ();
 FILLCELL_X2 FILLER_35_1 ();
 FILLCELL_X1 FILLER_35_3 ();
 FILLCELL_X2 FILLER_35_8 ();
 FILLCELL_X4 FILLER_35_14 ();
 FILLCELL_X2 FILLER_35_18 ();
 FILLCELL_X2 FILLER_35_23 ();
 FILLCELL_X2 FILLER_35_28 ();
 FILLCELL_X2 FILLER_35_33 ();
 FILLCELL_X2 FILLER_35_52 ();
 FILLCELL_X2 FILLER_35_58 ();
 FILLCELL_X4 FILLER_35_77 ();
 FILLCELL_X2 FILLER_35_81 ();
 FILLCELL_X2 FILLER_35_86 ();
 FILLCELL_X16 FILLER_35_92 ();
 FILLCELL_X2 FILLER_35_113 ();
 FILLCELL_X2 FILLER_35_124 ();
 FILLCELL_X16 FILLER_35_131 ();
 FILLCELL_X32 FILLER_35_148 ();
 FILLCELL_X32 FILLER_35_180 ();
 FILLCELL_X32 FILLER_35_212 ();
 FILLCELL_X32 FILLER_35_244 ();
 FILLCELL_X16 FILLER_35_276 ();
 FILLCELL_X2 FILLER_35_292 ();
 FILLCELL_X32 FILLER_35_295 ();
 FILLCELL_X32 FILLER_35_327 ();
 FILLCELL_X32 FILLER_35_359 ();
 FILLCELL_X16 FILLER_35_391 ();
 FILLCELL_X8 FILLER_35_407 ();
 FILLCELL_X4 FILLER_35_415 ();
 FILLCELL_X2 FILLER_35_419 ();
 FILLCELL_X4 FILLER_36_1 ();
 FILLCELL_X1 FILLER_36_5 ();
 FILLCELL_X2 FILLER_36_11 ();
 FILLCELL_X2 FILLER_36_18 ();
 FILLCELL_X2 FILLER_36_22 ();
 FILLCELL_X4 FILLER_36_28 ();
 FILLCELL_X2 FILLER_36_35 ();
 FILLCELL_X2 FILLER_36_42 ();
 FILLCELL_X2 FILLER_36_53 ();
 FILLCELL_X2 FILLER_36_58 ();
 FILLCELL_X2 FILLER_36_64 ();
 FILLCELL_X1 FILLER_36_66 ();
 FILLCELL_X2 FILLER_36_71 ();
 FILLCELL_X4 FILLER_36_74 ();
 FILLCELL_X1 FILLER_36_78 ();
 FILLCELL_X4 FILLER_36_86 ();
 FILLCELL_X2 FILLER_36_90 ();
 FILLCELL_X4 FILLER_36_109 ();
 FILLCELL_X32 FILLER_36_122 ();
 FILLCELL_X32 FILLER_36_154 ();
 FILLCELL_X32 FILLER_36_186 ();
 FILLCELL_X2 FILLER_36_218 ();
 FILLCELL_X32 FILLER_36_221 ();
 FILLCELL_X32 FILLER_36_253 ();
 FILLCELL_X32 FILLER_36_285 ();
 FILLCELL_X32 FILLER_36_317 ();
 FILLCELL_X16 FILLER_36_349 ();
 FILLCELL_X2 FILLER_36_365 ();
 FILLCELL_X32 FILLER_36_368 ();
 FILLCELL_X16 FILLER_36_400 ();
 FILLCELL_X4 FILLER_36_416 ();
 FILLCELL_X1 FILLER_36_420 ();
 FILLCELL_X4 FILLER_37_1 ();
 FILLCELL_X2 FILLER_37_8 ();
 FILLCELL_X4 FILLER_37_14 ();
 FILLCELL_X1 FILLER_37_18 ();
 FILLCELL_X2 FILLER_37_22 ();
 FILLCELL_X2 FILLER_37_27 ();
 FILLCELL_X2 FILLER_37_32 ();
 FILLCELL_X2 FILLER_37_44 ();
 FILLCELL_X2 FILLER_37_55 ();
 FILLCELL_X2 FILLER_37_66 ();
 FILLCELL_X2 FILLER_37_77 ();
 FILLCELL_X2 FILLER_37_92 ();
 FILLCELL_X2 FILLER_37_98 ();
 FILLCELL_X1 FILLER_37_100 ();
 FILLCELL_X2 FILLER_37_104 ();
 FILLCELL_X16 FILLER_37_119 ();
 FILLCELL_X8 FILLER_37_135 ();
 FILLCELL_X4 FILLER_37_143 ();
 FILLCELL_X32 FILLER_37_148 ();
 FILLCELL_X32 FILLER_37_180 ();
 FILLCELL_X32 FILLER_37_212 ();
 FILLCELL_X32 FILLER_37_244 ();
 FILLCELL_X16 FILLER_37_276 ();
 FILLCELL_X2 FILLER_37_292 ();
 FILLCELL_X32 FILLER_37_295 ();
 FILLCELL_X32 FILLER_37_327 ();
 FILLCELL_X32 FILLER_37_359 ();
 FILLCELL_X16 FILLER_37_391 ();
 FILLCELL_X8 FILLER_37_407 ();
 FILLCELL_X4 FILLER_37_415 ();
 FILLCELL_X2 FILLER_37_419 ();
 FILLCELL_X2 FILLER_38_1 ();
 FILLCELL_X2 FILLER_38_20 ();
 FILLCELL_X1 FILLER_38_22 ();
 FILLCELL_X2 FILLER_38_25 ();
 FILLCELL_X1 FILLER_38_27 ();
 FILLCELL_X2 FILLER_38_31 ();
 FILLCELL_X2 FILLER_38_43 ();
 FILLCELL_X2 FILLER_38_47 ();
 FILLCELL_X2 FILLER_38_59 ();
 FILLCELL_X2 FILLER_38_70 ();
 FILLCELL_X1 FILLER_38_72 ();
 FILLCELL_X2 FILLER_38_74 ();
 FILLCELL_X2 FILLER_38_94 ();
 FILLCELL_X4 FILLER_38_101 ();
 FILLCELL_X2 FILLER_38_105 ();
 FILLCELL_X32 FILLER_38_116 ();
 FILLCELL_X32 FILLER_38_148 ();
 FILLCELL_X32 FILLER_38_180 ();
 FILLCELL_X8 FILLER_38_212 ();
 FILLCELL_X32 FILLER_38_221 ();
 FILLCELL_X32 FILLER_38_253 ();
 FILLCELL_X32 FILLER_38_285 ();
 FILLCELL_X32 FILLER_38_317 ();
 FILLCELL_X16 FILLER_38_349 ();
 FILLCELL_X2 FILLER_38_365 ();
 FILLCELL_X32 FILLER_38_368 ();
 FILLCELL_X16 FILLER_38_400 ();
 FILLCELL_X4 FILLER_38_416 ();
 FILLCELL_X1 FILLER_38_420 ();
 FILLCELL_X4 FILLER_39_1 ();
 FILLCELL_X2 FILLER_39_22 ();
 FILLCELL_X8 FILLER_39_27 ();
 FILLCELL_X4 FILLER_39_35 ();
 FILLCELL_X1 FILLER_39_39 ();
 FILLCELL_X2 FILLER_39_44 ();
 FILLCELL_X2 FILLER_39_56 ();
 FILLCELL_X8 FILLER_39_67 ();
 FILLCELL_X4 FILLER_39_75 ();
 FILLCELL_X2 FILLER_39_79 ();
 FILLCELL_X1 FILLER_39_81 ();
 FILLCELL_X32 FILLER_39_91 ();
 FILLCELL_X16 FILLER_39_123 ();
 FILLCELL_X8 FILLER_39_139 ();
 FILLCELL_X32 FILLER_39_148 ();
 FILLCELL_X32 FILLER_39_180 ();
 FILLCELL_X32 FILLER_39_212 ();
 FILLCELL_X32 FILLER_39_244 ();
 FILLCELL_X16 FILLER_39_276 ();
 FILLCELL_X2 FILLER_39_292 ();
 FILLCELL_X32 FILLER_39_295 ();
 FILLCELL_X32 FILLER_39_327 ();
 FILLCELL_X32 FILLER_39_359 ();
 FILLCELL_X16 FILLER_39_391 ();
 FILLCELL_X8 FILLER_39_407 ();
 FILLCELL_X4 FILLER_39_415 ();
 FILLCELL_X2 FILLER_39_419 ();
 FILLCELL_X16 FILLER_40_1 ();
 FILLCELL_X1 FILLER_40_17 ();
 FILLCELL_X2 FILLER_40_35 ();
 FILLCELL_X1 FILLER_40_37 ();
 FILLCELL_X2 FILLER_40_55 ();
 FILLCELL_X8 FILLER_40_60 ();
 FILLCELL_X4 FILLER_40_68 ();
 FILLCELL_X1 FILLER_40_72 ();
 FILLCELL_X32 FILLER_40_74 ();
 FILLCELL_X32 FILLER_40_106 ();
 FILLCELL_X32 FILLER_40_138 ();
 FILLCELL_X32 FILLER_40_170 ();
 FILLCELL_X16 FILLER_40_202 ();
 FILLCELL_X2 FILLER_40_218 ();
 FILLCELL_X32 FILLER_40_221 ();
 FILLCELL_X32 FILLER_40_253 ();
 FILLCELL_X32 FILLER_40_285 ();
 FILLCELL_X32 FILLER_40_317 ();
 FILLCELL_X16 FILLER_40_349 ();
 FILLCELL_X2 FILLER_40_365 ();
 FILLCELL_X32 FILLER_40_368 ();
 FILLCELL_X16 FILLER_40_400 ();
 FILLCELL_X4 FILLER_40_416 ();
 FILLCELL_X1 FILLER_40_420 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X16 FILLER_41_33 ();
 FILLCELL_X4 FILLER_41_49 ();
 FILLCELL_X32 FILLER_41_55 ();
 FILLCELL_X32 FILLER_41_87 ();
 FILLCELL_X16 FILLER_41_119 ();
 FILLCELL_X8 FILLER_41_135 ();
 FILLCELL_X4 FILLER_41_143 ();
 FILLCELL_X32 FILLER_41_148 ();
 FILLCELL_X32 FILLER_41_180 ();
 FILLCELL_X32 FILLER_41_212 ();
 FILLCELL_X32 FILLER_41_244 ();
 FILLCELL_X16 FILLER_41_276 ();
 FILLCELL_X2 FILLER_41_292 ();
 FILLCELL_X32 FILLER_41_295 ();
 FILLCELL_X32 FILLER_41_327 ();
 FILLCELL_X32 FILLER_41_359 ();
 FILLCELL_X16 FILLER_41_391 ();
 FILLCELL_X8 FILLER_41_407 ();
 FILLCELL_X4 FILLER_41_415 ();
 FILLCELL_X2 FILLER_41_419 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X8 FILLER_42_65 ();
 FILLCELL_X32 FILLER_42_74 ();
 FILLCELL_X32 FILLER_42_106 ();
 FILLCELL_X32 FILLER_42_138 ();
 FILLCELL_X32 FILLER_42_170 ();
 FILLCELL_X16 FILLER_42_202 ();
 FILLCELL_X2 FILLER_42_218 ();
 FILLCELL_X32 FILLER_42_221 ();
 FILLCELL_X32 FILLER_42_253 ();
 FILLCELL_X32 FILLER_42_285 ();
 FILLCELL_X32 FILLER_42_317 ();
 FILLCELL_X16 FILLER_42_349 ();
 FILLCELL_X2 FILLER_42_365 ();
 FILLCELL_X32 FILLER_42_368 ();
 FILLCELL_X16 FILLER_42_400 ();
 FILLCELL_X4 FILLER_42_416 ();
 FILLCELL_X1 FILLER_42_420 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X32 FILLER_43_65 ();
 FILLCELL_X32 FILLER_43_97 ();
 FILLCELL_X16 FILLER_43_129 ();
 FILLCELL_X2 FILLER_43_145 ();
 FILLCELL_X32 FILLER_43_148 ();
 FILLCELL_X32 FILLER_43_180 ();
 FILLCELL_X32 FILLER_43_212 ();
 FILLCELL_X32 FILLER_43_244 ();
 FILLCELL_X16 FILLER_43_276 ();
 FILLCELL_X2 FILLER_43_292 ();
 FILLCELL_X32 FILLER_43_295 ();
 FILLCELL_X32 FILLER_43_327 ();
 FILLCELL_X32 FILLER_43_359 ();
 FILLCELL_X16 FILLER_43_391 ();
 FILLCELL_X8 FILLER_43_407 ();
 FILLCELL_X4 FILLER_43_415 ();
 FILLCELL_X2 FILLER_43_419 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X32 FILLER_44_33 ();
 FILLCELL_X8 FILLER_44_65 ();
 FILLCELL_X32 FILLER_44_74 ();
 FILLCELL_X32 FILLER_44_106 ();
 FILLCELL_X32 FILLER_44_138 ();
 FILLCELL_X32 FILLER_44_170 ();
 FILLCELL_X16 FILLER_44_202 ();
 FILLCELL_X2 FILLER_44_218 ();
 FILLCELL_X32 FILLER_44_221 ();
 FILLCELL_X32 FILLER_44_253 ();
 FILLCELL_X32 FILLER_44_285 ();
 FILLCELL_X32 FILLER_44_317 ();
 FILLCELL_X16 FILLER_44_349 ();
 FILLCELL_X2 FILLER_44_365 ();
 FILLCELL_X32 FILLER_44_368 ();
 FILLCELL_X16 FILLER_44_400 ();
 FILLCELL_X4 FILLER_44_416 ();
 FILLCELL_X1 FILLER_44_420 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X32 FILLER_45_33 ();
 FILLCELL_X32 FILLER_45_65 ();
 FILLCELL_X32 FILLER_45_97 ();
 FILLCELL_X16 FILLER_45_129 ();
 FILLCELL_X2 FILLER_45_145 ();
 FILLCELL_X32 FILLER_45_148 ();
 FILLCELL_X32 FILLER_45_180 ();
 FILLCELL_X32 FILLER_45_212 ();
 FILLCELL_X32 FILLER_45_244 ();
 FILLCELL_X16 FILLER_45_276 ();
 FILLCELL_X2 FILLER_45_292 ();
 FILLCELL_X32 FILLER_45_295 ();
 FILLCELL_X32 FILLER_45_327 ();
 FILLCELL_X32 FILLER_45_359 ();
 FILLCELL_X16 FILLER_45_391 ();
 FILLCELL_X8 FILLER_45_407 ();
 FILLCELL_X4 FILLER_45_415 ();
 FILLCELL_X2 FILLER_45_419 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X32 FILLER_46_33 ();
 FILLCELL_X8 FILLER_46_65 ();
 FILLCELL_X32 FILLER_46_74 ();
 FILLCELL_X32 FILLER_46_106 ();
 FILLCELL_X32 FILLER_46_138 ();
 FILLCELL_X32 FILLER_46_170 ();
 FILLCELL_X16 FILLER_46_202 ();
 FILLCELL_X2 FILLER_46_218 ();
 FILLCELL_X32 FILLER_46_221 ();
 FILLCELL_X32 FILLER_46_253 ();
 FILLCELL_X32 FILLER_46_285 ();
 FILLCELL_X32 FILLER_46_317 ();
 FILLCELL_X16 FILLER_46_349 ();
 FILLCELL_X2 FILLER_46_365 ();
 FILLCELL_X32 FILLER_46_368 ();
 FILLCELL_X16 FILLER_46_400 ();
 FILLCELL_X4 FILLER_46_416 ();
 FILLCELL_X1 FILLER_46_420 ();
 FILLCELL_X32 FILLER_47_1 ();
 FILLCELL_X32 FILLER_47_33 ();
 FILLCELL_X32 FILLER_47_65 ();
 FILLCELL_X32 FILLER_47_97 ();
 FILLCELL_X16 FILLER_47_129 ();
 FILLCELL_X2 FILLER_47_145 ();
 FILLCELL_X32 FILLER_47_148 ();
 FILLCELL_X32 FILLER_47_180 ();
 FILLCELL_X32 FILLER_47_212 ();
 FILLCELL_X32 FILLER_47_244 ();
 FILLCELL_X16 FILLER_47_276 ();
 FILLCELL_X2 FILLER_47_292 ();
 FILLCELL_X32 FILLER_47_295 ();
 FILLCELL_X32 FILLER_47_327 ();
 FILLCELL_X32 FILLER_47_359 ();
 FILLCELL_X16 FILLER_47_391 ();
 FILLCELL_X8 FILLER_47_407 ();
 FILLCELL_X4 FILLER_47_415 ();
 FILLCELL_X2 FILLER_47_419 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X32 FILLER_48_33 ();
 FILLCELL_X8 FILLER_48_65 ();
 FILLCELL_X32 FILLER_48_74 ();
 FILLCELL_X32 FILLER_48_106 ();
 FILLCELL_X32 FILLER_48_138 ();
 FILLCELL_X32 FILLER_48_170 ();
 FILLCELL_X16 FILLER_48_202 ();
 FILLCELL_X2 FILLER_48_218 ();
 FILLCELL_X32 FILLER_48_221 ();
 FILLCELL_X32 FILLER_48_253 ();
 FILLCELL_X32 FILLER_48_285 ();
 FILLCELL_X32 FILLER_48_317 ();
 FILLCELL_X16 FILLER_48_349 ();
 FILLCELL_X2 FILLER_48_365 ();
 FILLCELL_X32 FILLER_48_368 ();
 FILLCELL_X16 FILLER_48_400 ();
 FILLCELL_X4 FILLER_48_416 ();
 FILLCELL_X1 FILLER_48_420 ();
 FILLCELL_X32 FILLER_49_1 ();
 FILLCELL_X32 FILLER_49_33 ();
 FILLCELL_X32 FILLER_49_65 ();
 FILLCELL_X32 FILLER_49_97 ();
 FILLCELL_X16 FILLER_49_129 ();
 FILLCELL_X2 FILLER_49_145 ();
 FILLCELL_X32 FILLER_49_148 ();
 FILLCELL_X32 FILLER_49_180 ();
 FILLCELL_X32 FILLER_49_212 ();
 FILLCELL_X32 FILLER_49_244 ();
 FILLCELL_X16 FILLER_49_276 ();
 FILLCELL_X2 FILLER_49_292 ();
 FILLCELL_X32 FILLER_49_295 ();
 FILLCELL_X32 FILLER_49_327 ();
 FILLCELL_X32 FILLER_49_359 ();
 FILLCELL_X16 FILLER_49_391 ();
 FILLCELL_X8 FILLER_49_407 ();
 FILLCELL_X4 FILLER_49_415 ();
 FILLCELL_X2 FILLER_49_419 ();
 FILLCELL_X32 FILLER_50_1 ();
 FILLCELL_X32 FILLER_50_33 ();
 FILLCELL_X8 FILLER_50_65 ();
 FILLCELL_X32 FILLER_50_74 ();
 FILLCELL_X32 FILLER_50_106 ();
 FILLCELL_X32 FILLER_50_138 ();
 FILLCELL_X32 FILLER_50_170 ();
 FILLCELL_X16 FILLER_50_202 ();
 FILLCELL_X2 FILLER_50_218 ();
 FILLCELL_X32 FILLER_50_221 ();
 FILLCELL_X32 FILLER_50_253 ();
 FILLCELL_X32 FILLER_50_285 ();
 FILLCELL_X32 FILLER_50_317 ();
 FILLCELL_X16 FILLER_50_349 ();
 FILLCELL_X2 FILLER_50_365 ();
 FILLCELL_X32 FILLER_50_368 ();
 FILLCELL_X16 FILLER_50_400 ();
 FILLCELL_X4 FILLER_50_416 ();
 FILLCELL_X1 FILLER_50_420 ();
 FILLCELL_X32 FILLER_51_1 ();
 FILLCELL_X32 FILLER_51_33 ();
 FILLCELL_X32 FILLER_51_65 ();
 FILLCELL_X32 FILLER_51_97 ();
 FILLCELL_X16 FILLER_51_129 ();
 FILLCELL_X2 FILLER_51_145 ();
 FILLCELL_X32 FILLER_51_148 ();
 FILLCELL_X32 FILLER_51_180 ();
 FILLCELL_X32 FILLER_51_212 ();
 FILLCELL_X32 FILLER_51_244 ();
 FILLCELL_X16 FILLER_51_276 ();
 FILLCELL_X2 FILLER_51_292 ();
 FILLCELL_X32 FILLER_51_295 ();
 FILLCELL_X32 FILLER_51_327 ();
 FILLCELL_X32 FILLER_51_359 ();
 FILLCELL_X16 FILLER_51_391 ();
 FILLCELL_X8 FILLER_51_407 ();
 FILLCELL_X4 FILLER_51_415 ();
 FILLCELL_X2 FILLER_51_419 ();
 FILLCELL_X32 FILLER_52_1 ();
 FILLCELL_X32 FILLER_52_33 ();
 FILLCELL_X8 FILLER_52_65 ();
 FILLCELL_X32 FILLER_52_74 ();
 FILLCELL_X32 FILLER_52_106 ();
 FILLCELL_X32 FILLER_52_138 ();
 FILLCELL_X32 FILLER_52_170 ();
 FILLCELL_X16 FILLER_52_202 ();
 FILLCELL_X2 FILLER_52_218 ();
 FILLCELL_X32 FILLER_52_221 ();
 FILLCELL_X32 FILLER_52_253 ();
 FILLCELL_X32 FILLER_52_285 ();
 FILLCELL_X32 FILLER_52_317 ();
 FILLCELL_X16 FILLER_52_349 ();
 FILLCELL_X2 FILLER_52_365 ();
 FILLCELL_X32 FILLER_52_368 ();
 FILLCELL_X16 FILLER_52_400 ();
 FILLCELL_X4 FILLER_52_416 ();
 FILLCELL_X1 FILLER_52_420 ();
 FILLCELL_X32 FILLER_53_1 ();
 FILLCELL_X32 FILLER_53_33 ();
 FILLCELL_X32 FILLER_53_65 ();
 FILLCELL_X32 FILLER_53_97 ();
 FILLCELL_X16 FILLER_53_129 ();
 FILLCELL_X2 FILLER_53_145 ();
 FILLCELL_X32 FILLER_53_148 ();
 FILLCELL_X32 FILLER_53_180 ();
 FILLCELL_X32 FILLER_53_212 ();
 FILLCELL_X32 FILLER_53_244 ();
 FILLCELL_X16 FILLER_53_276 ();
 FILLCELL_X2 FILLER_53_292 ();
 FILLCELL_X32 FILLER_53_295 ();
 FILLCELL_X32 FILLER_53_327 ();
 FILLCELL_X32 FILLER_53_359 ();
 FILLCELL_X16 FILLER_53_391 ();
 FILLCELL_X8 FILLER_53_407 ();
 FILLCELL_X4 FILLER_53_415 ();
 FILLCELL_X2 FILLER_53_419 ();
 FILLCELL_X32 FILLER_54_1 ();
 FILLCELL_X32 FILLER_54_33 ();
 FILLCELL_X8 FILLER_54_65 ();
 FILLCELL_X32 FILLER_54_74 ();
 FILLCELL_X32 FILLER_54_106 ();
 FILLCELL_X32 FILLER_54_138 ();
 FILLCELL_X32 FILLER_54_170 ();
 FILLCELL_X16 FILLER_54_202 ();
 FILLCELL_X2 FILLER_54_218 ();
 FILLCELL_X32 FILLER_54_221 ();
 FILLCELL_X32 FILLER_54_253 ();
 FILLCELL_X32 FILLER_54_285 ();
 FILLCELL_X32 FILLER_54_317 ();
 FILLCELL_X16 FILLER_54_349 ();
 FILLCELL_X2 FILLER_54_365 ();
 FILLCELL_X32 FILLER_54_368 ();
 FILLCELL_X16 FILLER_54_400 ();
 FILLCELL_X4 FILLER_54_416 ();
 FILLCELL_X1 FILLER_54_420 ();
 FILLCELL_X32 FILLER_55_1 ();
 FILLCELL_X32 FILLER_55_33 ();
 FILLCELL_X32 FILLER_55_65 ();
 FILLCELL_X32 FILLER_55_97 ();
 FILLCELL_X16 FILLER_55_129 ();
 FILLCELL_X2 FILLER_55_145 ();
 FILLCELL_X32 FILLER_55_148 ();
 FILLCELL_X32 FILLER_55_180 ();
 FILLCELL_X32 FILLER_55_212 ();
 FILLCELL_X32 FILLER_55_244 ();
 FILLCELL_X16 FILLER_55_276 ();
 FILLCELL_X2 FILLER_55_292 ();
 FILLCELL_X32 FILLER_55_295 ();
 FILLCELL_X32 FILLER_55_327 ();
 FILLCELL_X32 FILLER_55_359 ();
 FILLCELL_X16 FILLER_55_391 ();
 FILLCELL_X8 FILLER_55_407 ();
 FILLCELL_X4 FILLER_55_415 ();
 FILLCELL_X2 FILLER_55_419 ();
 FILLCELL_X32 FILLER_56_1 ();
 FILLCELL_X32 FILLER_56_33 ();
 FILLCELL_X8 FILLER_56_65 ();
 FILLCELL_X32 FILLER_56_74 ();
 FILLCELL_X32 FILLER_56_106 ();
 FILLCELL_X8 FILLER_56_138 ();
 FILLCELL_X32 FILLER_56_147 ();
 FILLCELL_X32 FILLER_56_179 ();
 FILLCELL_X8 FILLER_56_211 ();
 FILLCELL_X32 FILLER_56_220 ();
 FILLCELL_X32 FILLER_56_252 ();
 FILLCELL_X8 FILLER_56_284 ();
 FILLCELL_X32 FILLER_56_293 ();
 FILLCELL_X32 FILLER_56_325 ();
 FILLCELL_X8 FILLER_56_357 ();
 FILLCELL_X32 FILLER_56_366 ();
 FILLCELL_X16 FILLER_56_398 ();
 FILLCELL_X4 FILLER_56_414 ();
 FILLCELL_X2 FILLER_56_418 ();
 FILLCELL_X1 FILLER_56_420 ();
endmodule
